// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 14.1.1 Build 190 01/19/2015 SJ Web Edition"

// DATE "05/06/2015 19:06:06"

// 
// Device: Altera EP4CE115F29C7 Package FBGA780
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module usb_system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	all_switches_wire_export,
	clk_clk,
	keycode_export,
	led_wire_export,
	red_leds_wire_export,
	reset_reset_n,
	sdram_out_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	usb_DATA,
	usb_ADDR,
	usb_RD_N,
	usb_WR_N,
	usb_CS_N,
	usb_RST_N,
	usb_INT,
	usb_out_clk_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	[17:0] all_switches_wire_export;
input 	clk_clk;
output 	[7:0] keycode_export;
output 	[7:0] led_wire_export;
output 	[17:0] red_leds_wire_export;
input 	reset_reset_n;
output 	sdram_out_clk_clk;
output 	[12:0] sdram_wire_addr;
output 	[1:0] sdram_wire_ba;
output 	sdram_wire_cas_n;
output 	sdram_wire_cke;
output 	sdram_wire_cs_n;
inout 	[31:0] sdram_wire_dq;
output 	[3:0] sdram_wire_dqm;
output 	sdram_wire_ras_n;
output 	sdram_wire_we_n;
inout 	[15:0] usb_DATA;
output 	[1:0] usb_ADDR;
output 	usb_RD_N;
output 	usb_WR_N;
output 	usb_CS_N;
output 	usb_RST_N;
input 	usb_INT;
output 	usb_out_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clocks|sd1|wire_pll7_clk[0] ;
wire \clocks|sd1|wire_pll7_clk[1] ;
wire \sdram|m_addr[0]~q ;
wire \sdram|m_addr[1]~q ;
wire \sdram|m_addr[2]~q ;
wire \sdram|m_addr[3]~q ;
wire \sdram|m_addr[4]~q ;
wire \sdram|m_addr[5]~q ;
wire \sdram|m_addr[6]~q ;
wire \sdram|m_addr[7]~q ;
wire \sdram|m_addr[8]~q ;
wire \sdram|m_addr[9]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|sr[0]~q ;
wire \cpu|cpu|W_alu_result[7]~q ;
wire \cpu|cpu|W_alu_result[14]~q ;
wire \cpu|cpu|W_alu_result[13]~q ;
wire \cpu|cpu|W_alu_result[18]~q ;
wire \cpu|cpu|W_alu_result[17]~q ;
wire \cpu|cpu|W_alu_result[16]~q ;
wire \cpu|cpu|W_alu_result[15]~q ;
wire \cpu|cpu|W_alu_result[12]~q ;
wire \cpu|cpu|W_alu_result[11]~q ;
wire \cpu|cpu|W_alu_result[10]~q ;
wire \cpu|cpu|W_alu_result[9]~q ;
wire \cpu|cpu|W_alu_result[23]~q ;
wire \cpu|cpu|W_alu_result[22]~q ;
wire \cpu|cpu|W_alu_result[8]~q ;
wire \cpu|cpu|W_alu_result[6]~q ;
wire \cpu|cpu|W_alu_result[24]~q ;
wire \cpu|cpu|W_alu_result[21]~q ;
wire \cpu|cpu|W_alu_result[20]~q ;
wire \cpu|cpu|W_alu_result[19]~q ;
wire \cpu|cpu|W_alu_result[28]~q ;
wire \cpu|cpu|W_alu_result[27]~q ;
wire \cpu|cpu|W_alu_result[26]~q ;
wire \cpu|cpu|W_alu_result[25]~q ;
wire \cpu|cpu|W_alu_result[4]~q ;
wire \cpu|cpu|W_alu_result[5]~q ;
wire \cpu|cpu|W_alu_result[2]~q ;
wire \cpu|cpu|W_alu_result[3]~q ;
wire \sdram|oe~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[0]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[1]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[2]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[3]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[5]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[6]~q ;
wire \cpu|cpu|d_writedata[24]~q ;
wire \cpu|cpu|d_writedata[25]~q ;
wire \cpu|cpu|d_writedata[26]~q ;
wire \cpu|cpu|d_writedata[27]~q ;
wire \cpu|cpu|d_writedata[28]~q ;
wire \cpu|cpu|d_writedata[29]~q ;
wire \cpu|cpu|d_writedata[30]~q ;
wire \cpu|cpu|d_writedata[31]~q ;
wire \keycode|data_out[0]~q ;
wire \keycode|data_out[1]~q ;
wire \keycode|data_out[2]~q ;
wire \keycode|data_out[3]~q ;
wire \keycode|data_out[4]~q ;
wire \keycode|data_out[5]~q ;
wire \keycode|data_out[6]~q ;
wire \keycode|data_out[7]~q ;
wire \led|data_out[0]~q ;
wire \led|data_out[1]~q ;
wire \led|data_out[2]~q ;
wire \led|data_out[3]~q ;
wire \led|data_out[4]~q ;
wire \led|data_out[5]~q ;
wire \led|data_out[6]~q ;
wire \led|data_out[7]~q ;
wire \red_leds|data_out[0]~q ;
wire \red_leds|data_out[1]~q ;
wire \red_leds|data_out[2]~q ;
wire \red_leds|data_out[3]~q ;
wire \red_leds|data_out[4]~q ;
wire \red_leds|data_out[5]~q ;
wire \red_leds|data_out[6]~q ;
wire \red_leds|data_out[7]~q ;
wire \red_leds|data_out[8]~q ;
wire \red_leds|data_out[9]~q ;
wire \red_leds|data_out[10]~q ;
wire \red_leds|data_out[11]~q ;
wire \red_leds|data_out[12]~q ;
wire \red_leds|data_out[13]~q ;
wire \red_leds|data_out[14]~q ;
wire \red_leds|data_out[15]~q ;
wire \red_leds|data_out[16]~q ;
wire \red_leds|data_out[17]~q ;
wire \sdram|m_addr[10]~q ;
wire \sdram|m_addr[11]~q ;
wire \sdram|m_addr[12]~q ;
wire \sdram|m_bank[0]~q ;
wire \sdram|m_bank[1]~q ;
wire \sdram|m_cmd[1]~q ;
wire \sdram|m_cmd[3]~q ;
wire \sdram|m_dqm[0]~q ;
wire \sdram|m_dqm[1]~q ;
wire \sdram|m_dqm[2]~q ;
wire \sdram|m_dqm[3]~q ;
wire \sdram|m_cmd[2]~q ;
wire \sdram|m_cmd[0]~q ;
wire \cy7c67200_if_0|HPI_ADDR[0]~q ;
wire \cy7c67200_if_0|HPI_ADDR[1]~q ;
wire \cy7c67200_if_0|HPI_RD_N~q ;
wire \cy7c67200_if_0|HPI_WR_N~q ;
wire \cy7c67200_if_0|HPI_CS_N~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|ir_out[0]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|ir_out[1]~q ;
wire \jtag_uart|usb_system_jtag_uart_alt_jtag_atlantic|tdo~q ;
wire \cpu|cpu|d_writedata[0]~q ;
wire \rst_controller_002|r_sync_rst~q ;
wire \mm_interconnect_0|router|Equal3~4_combout ;
wire \mm_interconnect_0|router|Equal6~0_combout ;
wire \mm_interconnect_0|keycode_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \keycode|always0~0_combout ;
wire \cpu|cpu|d_write~q ;
wire \mm_interconnect_0|cpu_data_master_translator|write_accepted~q ;
wire \keycode|always0~1_combout ;
wire \mm_interconnect_0|keycode_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|keycode_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|cpu|d_writedata[1]~q ;
wire \cpu|cpu|d_writedata[2]~q ;
wire \cpu|cpu|d_writedata[3]~q ;
wire \cpu|cpu|d_writedata[4]~q ;
wire \cpu|cpu|d_writedata[5]~q ;
wire \cpu|cpu|d_writedata[6]~q ;
wire \cpu|cpu|d_writedata[7]~q ;
wire \rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \led|always0~1_combout ;
wire \mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|red_leds_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \red_leds|always0~1_combout ;
wire \mm_interconnect_0|red_leds_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|red_leds_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|cpu|d_writedata[8]~q ;
wire \cpu|cpu|d_writedata[9]~q ;
wire \cpu|cpu|d_writedata[10]~q ;
wire \cpu|cpu|d_writedata[11]~q ;
wire \cpu|cpu|d_writedata[12]~q ;
wire \cpu|cpu|d_writedata[13]~q ;
wire \cpu|cpu|d_writedata[14]~q ;
wire \cpu|cpu|d_writedata[15]~q ;
wire \cpu|cpu|d_writedata[16]~q ;
wire \cpu|cpu|d_writedata[17]~q ;
wire \sdram|the_usb_system_sdram_input_efifo_module|entries[1]~q ;
wire \sdram|the_usb_system_sdram_input_efifo_module|entries[0]~q ;
wire \rst_controller_003|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[42]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[43]~q ;
wire \clock_crossing_io|cmd_fifo|out_valid~q ;
wire \clock_crossing_io|m0_read~0_combout ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_read~0_combout ;
wire \clock_crossing_io|cmd_fifo|out_payload[37]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_write~0_combout ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_oci_debug|resetrequest~q ;
wire \rst_controller|merged_reset~0_combout ;
wire \clock_crossing_io|cmd_fifo|sink_in_reset~q ;
wire \cpu|cpu|d_read~q ;
wire \mm_interconnect_0|cpu_data_master_translator|read_accepted~q ;
wire \mm_interconnect_0|keycode_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|red_leds_s1_translator|read_latency_shift_reg[0]~q ;
wire \clock_crossing_io|rsp_fifo|out_valid~q ;
wire \mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ;
wire \mm_interconnect_0|led_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|all_switches_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|clock_crossing_io_s0_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ;
wire \mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|keycode_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|led_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|red_leds_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|all_switches_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[67]~q ;
wire \cpu|cpu|av_ld_getting_data~6_combout ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ;
wire \mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \clock_crossing_io|cmd_fifo|full~q ;
wire \cpu|cpu|F_pc[26]~q ;
wire \cpu|cpu|F_pc[25]~q ;
wire \cpu|cpu|F_pc[24]~q ;
wire \cpu|cpu|F_pc[23]~q ;
wire \cpu|cpu|F_pc[22]~q ;
wire \cpu|cpu|F_pc[21]~q ;
wire \cpu|cpu|F_pc[20]~q ;
wire \cpu|cpu|F_pc[19]~q ;
wire \cpu|cpu|F_pc[18]~q ;
wire \cpu|cpu|F_pc[17]~q ;
wire \cpu|cpu|F_pc[16]~q ;
wire \cpu|cpu|F_pc[15]~q ;
wire \cpu|cpu|F_pc[14]~q ;
wire \cpu|cpu|F_pc[13]~q ;
wire \cpu|cpu|F_pc[12]~q ;
wire \cpu|cpu|F_pc[11]~q ;
wire \cpu|cpu|F_pc[10]~q ;
wire \cpu|cpu|F_pc[9]~q ;
wire \cpu|cpu|F_pc[8]~q ;
wire \cpu|cpu|F_pc[7]~q ;
wire \cpu|cpu|F_pc[5]~q ;
wire \cpu|cpu|F_pc[6]~q ;
wire \cpu|cpu|F_pc[4]~q ;
wire \cpu|cpu|F_pc[1]~q ;
wire \cpu|cpu|F_pc[3]~q ;
wire \cpu|cpu|i_read~q ;
wire \cpu|cpu|F_pc[2]~q ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \jtag_uart|av_waitrequest~q ;
wire \mm_interconnect_0|router|Equal9~1_combout ;
wire \mm_interconnect_0|cpu_data_master_translator|av_waitrequest~1_combout ;
wire \clock_crossing_io|s0_cmd_valid~combout ;
wire \mm_interconnect_0|cmd_mux_003|WideOr1~combout ;
wire \cpu|cpu|F_pc[0]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[38]~combout ;
wire \mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem~0_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_006|last_cycle~0_combout ;
wire \mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ;
wire \mm_interconnect_0|cmd_mux_006|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[68]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[62]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[51]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[50]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[53]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[52]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[55]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[54]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[57]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[56]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[59]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[58]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[61]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[60]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[47]~combout ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[32]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[32]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[33]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[33]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[34]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[34]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[35]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[35]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|waitrequest_reset_override~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_waitrequest_generated~1_combout ;
wire \sdram|m_data[0]~q ;
wire \sdram|m_data[1]~q ;
wire \sdram|m_data[2]~q ;
wire \sdram|m_data[3]~q ;
wire \sdram|m_data[4]~q ;
wire \sdram|m_data[5]~q ;
wire \sdram|m_data[6]~q ;
wire \sdram|m_data[7]~q ;
wire \sdram|m_data[8]~q ;
wire \sdram|m_data[9]~q ;
wire \sdram|m_data[10]~q ;
wire \sdram|m_data[11]~q ;
wire \sdram|m_data[12]~q ;
wire \sdram|m_data[13]~q ;
wire \sdram|m_data[14]~q ;
wire \sdram|m_data[15]~q ;
wire \sdram|m_data[16]~q ;
wire \sdram|m_data[17]~q ;
wire \sdram|m_data[18]~q ;
wire \sdram|m_data[19]~q ;
wire \sdram|m_data[20]~q ;
wire \sdram|m_data[21]~q ;
wire \sdram|m_data[22]~q ;
wire \sdram|m_data[23]~q ;
wire \sdram|m_data[24]~q ;
wire \sdram|m_data[25]~q ;
wire \sdram|m_data[26]~q ;
wire \sdram|m_data[27]~q ;
wire \sdram|m_data[28]~q ;
wire \sdram|m_data[29]~q ;
wire \sdram|m_data[30]~q ;
wire \sdram|m_data[31]~q ;
wire \cy7c67200_if_0|TMP_DATA[0]~q ;
wire \cy7c67200_if_0|TMP_DATA[1]~q ;
wire \cy7c67200_if_0|TMP_DATA[2]~q ;
wire \cy7c67200_if_0|TMP_DATA[3]~q ;
wire \cy7c67200_if_0|TMP_DATA[4]~q ;
wire \cy7c67200_if_0|TMP_DATA[5]~q ;
wire \cy7c67200_if_0|TMP_DATA[6]~q ;
wire \cy7c67200_if_0|TMP_DATA[7]~q ;
wire \cy7c67200_if_0|TMP_DATA[8]~q ;
wire \cy7c67200_if_0|TMP_DATA[9]~q ;
wire \cy7c67200_if_0|TMP_DATA[10]~q ;
wire \cy7c67200_if_0|TMP_DATA[11]~q ;
wire \cy7c67200_if_0|TMP_DATA[12]~q ;
wire \cy7c67200_if_0|TMP_DATA[13]~q ;
wire \cy7c67200_if_0|TMP_DATA[14]~q ;
wire \cy7c67200_if_0|TMP_DATA[15]~q ;
wire \mm_interconnect_0|cmd_demux|sink_ready~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|WideOr1~combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent|local_read~0_combout ;
wire \mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem~1_combout ;
wire \mm_interconnect_0|clock_crossing_io_s0_agent|m0_write~2_combout ;
wire \mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ;
wire \mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~0_combout ;
wire \mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~1_combout ;
wire \mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~2_combout ;
wire \cpu|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[0]~q ;
wire \mm_interconnect_0|clocks_pll_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[1]~q ;
wire \mm_interconnect_0|clocks_pll_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[2]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[4]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|read_latency_shift_reg[0]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[5]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[6]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[7]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[8]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[9]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[10]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[11]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[12]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[13]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[14]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[15]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[16]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[17]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[18]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[19]~q ;
wire \clock_crossing_io|cmd_fifo|out_payload[20]~q ;
wire \clock_crossing_io|rsp_fifo|out_payload[0]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[22]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[23]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[24]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[26]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[11]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[13]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~3_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[12]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[5]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[14]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[15]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[10]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[9]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[8]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[7]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[6]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[18]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[19]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[17]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[27]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[28]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[31]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem~4_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[1]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~0_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[2]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~28_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~30_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[3]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~34_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[4]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~37_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[5]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~41_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[6]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~45_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[7]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~49_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[8]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~combout ;
wire \irq_synchronizer|sync|sync[0].u|dreg[1]~q ;
wire \jtag_uart|av_readdata[9]~combout ;
wire \jtag_uart|av_readdata[8]~0_combout ;
wire \clocks|readdata[0]~1_combout ;
wire \clocks|readdata[1]~2_combout ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[4]~q ;
wire \clock_crossing_io|rsp_fifo|out_payload[9]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[10]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[10]~59_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[11]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[12]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[12]~66_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[13]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[14]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[14]~72_combout ;
wire \clock_crossing_io|rsp_fifo|out_payload[15]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[16]~78_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[17]~combout ;
wire \cpu|cpu|d_byteenable[0]~q ;
wire \cpu|cpu|d_byteenable[1]~q ;
wire \cpu|cpu|d_byteenable[2]~q ;
wire \cpu|cpu|d_byteenable[3]~q ;
wire \rst_controller_002|r_early_rst~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~32_combout ;
wire \jtag_uart|read_0~q ;
wire \jtag_uart|av_readdata[0]~1_combout ;
wire \led|readdata[0]~combout ;
wire \keycode|readdata[0]~combout ;
wire \all_switches|readdata[0]~q ;
wire \red_leds|readdata[0]~combout ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[22]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[23]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[24]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[25]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[26]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[11]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[13]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[16]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[12]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[14]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[15]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[10]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[9]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[8]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[7]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[20]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[18]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[19]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[17]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~11_combout ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[21]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~12_combout ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[27]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~14_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~16_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~18_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~20_combout ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[24]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[28]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[28]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[27]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[31]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[26]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[30]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[25]~q ;
wire \cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[29]~q ;
wire \jtag_uart|av_readdata[1]~2_combout ;
wire \led|readdata[1]~combout ;
wire \keycode|readdata[1]~combout ;
wire \all_switches|readdata[1]~q ;
wire \red_leds|readdata[1]~combout ;
wire \jtag_uart|av_readdata[2]~3_combout ;
wire \led|readdata[2]~combout ;
wire \keycode|readdata[2]~combout ;
wire \all_switches|readdata[2]~q ;
wire \red_leds|readdata[2]~combout ;
wire \all_switches|readdata[3]~q ;
wire \red_leds|readdata[3]~combout ;
wire \jtag_uart|av_readdata[3]~4_combout ;
wire \led|readdata[3]~combout ;
wire \keycode|readdata[3]~combout ;
wire \jtag_uart|av_readdata[4]~5_combout ;
wire \led|readdata[4]~combout ;
wire \keycode|readdata[4]~combout ;
wire \all_switches|readdata[4]~q ;
wire \red_leds|readdata[4]~combout ;
wire \jtag_uart|av_readdata[5]~6_combout ;
wire \led|readdata[5]~combout ;
wire \keycode|readdata[5]~combout ;
wire \all_switches|readdata[5]~q ;
wire \red_leds|readdata[5]~combout ;
wire \jtag_uart|av_readdata[6]~7_combout ;
wire \led|readdata[6]~combout ;
wire \keycode|readdata[6]~combout ;
wire \all_switches|readdata[6]~q ;
wire \red_leds|readdata[6]~combout ;
wire \jtag_uart|av_readdata[7]~8_combout ;
wire \led|readdata[7]~combout ;
wire \keycode|readdata[7]~combout ;
wire \all_switches|readdata[7]~q ;
wire \red_leds|readdata[7]~combout ;
wire \all_switches|readdata[8]~q ;
wire \red_leds|readdata[8]~combout ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \all_switches|readdata[9]~q ;
wire \red_leds|readdata[9]~combout ;
wire \jtag_uart|ac~q ;
wire \all_switches|readdata[10]~q ;
wire \red_leds|readdata[10]~combout ;
wire \all_switches|readdata[11]~q ;
wire \red_leds|readdata[11]~combout ;
wire \all_switches|readdata[12]~q ;
wire \red_leds|readdata[12]~combout ;
wire \all_switches|readdata[13]~q ;
wire \red_leds|readdata[13]~combout ;
wire \jtag_uart|woverflow~q ;
wire \all_switches|readdata[14]~q ;
wire \red_leds|readdata[14]~combout ;
wire \all_switches|readdata[15]~q ;
wire \red_leds|readdata[15]~combout ;
wire \jtag_uart|rvalid~q ;
wire \all_switches|readdata[16]~q ;
wire \red_leds|readdata[16]~combout ;
wire \all_switches|readdata[17]~q ;
wire \red_leds|readdata[17]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[31]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[15]~q ;
wire \sdram|za_valid~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \cpu|cpu|d_writedata[18]~q ;
wire \cpu|cpu|d_writedata[19]~q ;
wire \cpu|cpu|d_writedata[20]~q ;
wire \cpu|cpu|d_writedata[21]~q ;
wire \cpu|cpu|d_writedata[22]~q ;
wire \cpu|cpu|d_writedata[23]~q ;
wire \cy7c67200_if_0|oDATA[0]~q ;
wire \cy7c67200_if_0|oDATA[1]~q ;
wire \cy7c67200_if_0|oDATA[2]~q ;
wire \cy7c67200_if_0|oDATA[3]~q ;
wire \cy7c67200_if_0|oDATA[4]~q ;
wire \cy7c67200_if_0|oDATA[5]~q ;
wire \cy7c67200_if_0|oDATA[6]~q ;
wire \cy7c67200_if_0|oDATA[7]~q ;
wire \cy7c67200_if_0|oDATA[8]~q ;
wire \cy7c67200_if_0|oINT~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \cy7c67200_if_0|oDATA[9]~q ;
wire \cy7c67200_if_0|oDATA[10]~q ;
wire \cy7c67200_if_0|oDATA[11]~q ;
wire \cy7c67200_if_0|oDATA[12]~q ;
wire \cy7c67200_if_0|oDATA[13]~q ;
wire \cy7c67200_if_0|oDATA[14]~q ;
wire \cy7c67200_if_0|oDATA[15]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~32_combout ;
wire \sdram|za_data[0]~q ;
wire \sdram|za_data[1]~q ;
wire \sdram|za_data[2]~q ;
wire \sdram|za_data[3]~q ;
wire \sdram|za_data[4]~q ;
wire \sdram|za_data[22]~q ;
wire \sdram|za_data[23]~q ;
wire \sdram|za_data[24]~q ;
wire \sdram|za_data[25]~q ;
wire \sdram|za_data[26]~q ;
wire \sdram|za_data[11]~q ;
wire \sdram|za_data[13]~q ;
wire \sdram|za_data[16]~q ;
wire \sdram|za_data[12]~q ;
wire \sdram|za_data[5]~q ;
wire \sdram|za_data[14]~q ;
wire \sdram|za_data[15]~q ;
wire \sdram|za_data[10]~q ;
wire \sdram|za_data[9]~q ;
wire \sdram|za_data[8]~q ;
wire \sdram|za_data[7]~q ;
wire \sdram|za_data[6]~q ;
wire \sdram|za_data[20]~q ;
wire \sdram|za_data[18]~q ;
wire \sdram|za_data[19]~q ;
wire \sdram|za_data[17]~q ;
wire \sdram|za_data[21]~q ;
wire \sdram|za_data[27]~q ;
wire \sdram|za_data[28]~q ;
wire \sdram|za_data[31]~q ;
wire \sdram|za_data[30]~q ;
wire \sdram|za_data[29]~q ;
wire \mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_begintransfer~2_combout ;
wire \mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ;
wire \mm_interconnect_0|clock_crossing_io_s0_agent|m0_read~2_combout ;
wire \mm_interconnect_0|clock_crossing_io_s0_agent|m0_write~3_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~84_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~85_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~86_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~87_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~88_combout ;
wire \rst_controller_002|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \sdram_wire_dq[0]~input_o ;
wire \sdram_wire_dq[1]~input_o ;
wire \sdram_wire_dq[2]~input_o ;
wire \sdram_wire_dq[3]~input_o ;
wire \sdram_wire_dq[4]~input_o ;
wire \sdram_wire_dq[5]~input_o ;
wire \sdram_wire_dq[6]~input_o ;
wire \sdram_wire_dq[7]~input_o ;
wire \sdram_wire_dq[8]~input_o ;
wire \sdram_wire_dq[9]~input_o ;
wire \sdram_wire_dq[10]~input_o ;
wire \sdram_wire_dq[11]~input_o ;
wire \sdram_wire_dq[12]~input_o ;
wire \sdram_wire_dq[13]~input_o ;
wire \sdram_wire_dq[14]~input_o ;
wire \sdram_wire_dq[15]~input_o ;
wire \sdram_wire_dq[16]~input_o ;
wire \sdram_wire_dq[17]~input_o ;
wire \sdram_wire_dq[18]~input_o ;
wire \sdram_wire_dq[19]~input_o ;
wire \sdram_wire_dq[20]~input_o ;
wire \sdram_wire_dq[21]~input_o ;
wire \sdram_wire_dq[22]~input_o ;
wire \sdram_wire_dq[23]~input_o ;
wire \sdram_wire_dq[24]~input_o ;
wire \sdram_wire_dq[25]~input_o ;
wire \sdram_wire_dq[26]~input_o ;
wire \sdram_wire_dq[27]~input_o ;
wire \sdram_wire_dq[28]~input_o ;
wire \sdram_wire_dq[29]~input_o ;
wire \sdram_wire_dq[30]~input_o ;
wire \sdram_wire_dq[31]~input_o ;
wire \usb_DATA[0]~input_o ;
wire \usb_DATA[1]~input_o ;
wire \usb_DATA[2]~input_o ;
wire \usb_DATA[3]~input_o ;
wire \usb_DATA[4]~input_o ;
wire \usb_DATA[5]~input_o ;
wire \usb_DATA[6]~input_o ;
wire \usb_DATA[7]~input_o ;
wire \usb_DATA[8]~input_o ;
wire \usb_DATA[9]~input_o ;
wire \usb_DATA[10]~input_o ;
wire \usb_DATA[11]~input_o ;
wire \usb_DATA[12]~input_o ;
wire \usb_DATA[13]~input_o ;
wire \usb_DATA[14]~input_o ;
wire \usb_DATA[15]~input_o ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \all_switches_wire_export[0]~input_o ;
wire \all_switches_wire_export[1]~input_o ;
wire \all_switches_wire_export[2]~input_o ;
wire \all_switches_wire_export[3]~input_o ;
wire \all_switches_wire_export[4]~input_o ;
wire \all_switches_wire_export[5]~input_o ;
wire \all_switches_wire_export[6]~input_o ;
wire \all_switches_wire_export[7]~input_o ;
wire \all_switches_wire_export[8]~input_o ;
wire \all_switches_wire_export[9]~input_o ;
wire \all_switches_wire_export[10]~input_o ;
wire \all_switches_wire_export[11]~input_o ;
wire \all_switches_wire_export[12]~input_o ;
wire \all_switches_wire_export[13]~input_o ;
wire \all_switches_wire_export[14]~input_o ;
wire \all_switches_wire_export[15]~input_o ;
wire \all_switches_wire_export[16]~input_o ;
wire \all_switches_wire_export[17]~input_o ;
wire \usb_INT~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~10 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;


usb_system_CY7C67200_IF cy7c67200_if_0(
	.iCLK(\clocks|sd1|wire_pll7_clk[1] ),
	.HPI_ADDR_0(\cy7c67200_if_0|HPI_ADDR[0]~q ),
	.HPI_ADDR_1(\cy7c67200_if_0|HPI_ADDR[1]~q ),
	.HPI_RD_N1(\cy7c67200_if_0|HPI_RD_N~q ),
	.HPI_WR_N1(\cy7c67200_if_0|HPI_WR_N~q ),
	.HPI_CS_N1(\cy7c67200_if_0|HPI_CS_N~q ),
	.iRST_N(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_payload_42(\clock_crossing_io|cmd_fifo|out_payload[42]~q ),
	.out_payload_43(\clock_crossing_io|cmd_fifo|out_payload[43]~q ),
	.av_read(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_read~0_combout ),
	.av_write(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_write~0_combout ),
	.TMP_DATA_0(\cy7c67200_if_0|TMP_DATA[0]~q ),
	.TMP_DATA_1(\cy7c67200_if_0|TMP_DATA[1]~q ),
	.TMP_DATA_2(\cy7c67200_if_0|TMP_DATA[2]~q ),
	.TMP_DATA_3(\cy7c67200_if_0|TMP_DATA[3]~q ),
	.TMP_DATA_4(\cy7c67200_if_0|TMP_DATA[4]~q ),
	.TMP_DATA_5(\cy7c67200_if_0|TMP_DATA[5]~q ),
	.TMP_DATA_6(\cy7c67200_if_0|TMP_DATA[6]~q ),
	.TMP_DATA_7(\cy7c67200_if_0|TMP_DATA[7]~q ),
	.TMP_DATA_8(\cy7c67200_if_0|TMP_DATA[8]~q ),
	.TMP_DATA_9(\cy7c67200_if_0|TMP_DATA[9]~q ),
	.TMP_DATA_10(\cy7c67200_if_0|TMP_DATA[10]~q ),
	.TMP_DATA_11(\cy7c67200_if_0|TMP_DATA[11]~q ),
	.TMP_DATA_12(\cy7c67200_if_0|TMP_DATA[12]~q ),
	.TMP_DATA_13(\cy7c67200_if_0|TMP_DATA[13]~q ),
	.TMP_DATA_14(\cy7c67200_if_0|TMP_DATA[14]~q ),
	.TMP_DATA_15(\cy7c67200_if_0|TMP_DATA[15]~q ),
	.iDATA({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\clock_crossing_io|cmd_fifo|out_payload[20]~q ,\clock_crossing_io|cmd_fifo|out_payload[19]~q ,\clock_crossing_io|cmd_fifo|out_payload[18]~q ,\clock_crossing_io|cmd_fifo|out_payload[17]~q ,
\clock_crossing_io|cmd_fifo|out_payload[16]~q ,\clock_crossing_io|cmd_fifo|out_payload[15]~q ,\clock_crossing_io|cmd_fifo|out_payload[14]~q ,\clock_crossing_io|cmd_fifo|out_payload[13]~q ,\clock_crossing_io|cmd_fifo|out_payload[12]~q ,
\clock_crossing_io|cmd_fifo|out_payload[11]~q ,\clock_crossing_io|cmd_fifo|out_payload[10]~q ,\clock_crossing_io|cmd_fifo|out_payload[9]~q ,\clock_crossing_io|cmd_fifo|out_payload[8]~q ,\clock_crossing_io|cmd_fifo|out_payload[7]~q ,
\clock_crossing_io|cmd_fifo|out_payload[6]~q ,\clock_crossing_io|cmd_fifo|out_payload[5]~q }),
	.oDATA_0(\cy7c67200_if_0|oDATA[0]~q ),
	.oDATA_1(\cy7c67200_if_0|oDATA[1]~q ),
	.oDATA_2(\cy7c67200_if_0|oDATA[2]~q ),
	.oDATA_3(\cy7c67200_if_0|oDATA[3]~q ),
	.oDATA_4(\cy7c67200_if_0|oDATA[4]~q ),
	.oDATA_5(\cy7c67200_if_0|oDATA[5]~q ),
	.oDATA_6(\cy7c67200_if_0|oDATA[6]~q ),
	.oDATA_7(\cy7c67200_if_0|oDATA[7]~q ),
	.oDATA_8(\cy7c67200_if_0|oDATA[8]~q ),
	.oINT1(\cy7c67200_if_0|oINT~q ),
	.oDATA_9(\cy7c67200_if_0|oDATA[9]~q ),
	.oDATA_10(\cy7c67200_if_0|oDATA[10]~q ),
	.oDATA_11(\cy7c67200_if_0|oDATA[11]~q ),
	.oDATA_12(\cy7c67200_if_0|oDATA[12]~q ),
	.oDATA_13(\cy7c67200_if_0|oDATA[13]~q ),
	.oDATA_14(\cy7c67200_if_0|oDATA[14]~q ),
	.oDATA_15(\cy7c67200_if_0|oDATA[15]~q ),
	.av_begintransfer(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_begintransfer~2_combout ),
	.usb_DATA_0(\usb_DATA[0]~input_o ),
	.usb_DATA_1(\usb_DATA[1]~input_o ),
	.usb_DATA_2(\usb_DATA[2]~input_o ),
	.usb_DATA_3(\usb_DATA[3]~input_o ),
	.usb_DATA_4(\usb_DATA[4]~input_o ),
	.usb_DATA_5(\usb_DATA[5]~input_o ),
	.usb_DATA_6(\usb_DATA[6]~input_o ),
	.usb_DATA_7(\usb_DATA[7]~input_o ),
	.usb_DATA_8(\usb_DATA[8]~input_o ),
	.usb_DATA_9(\usb_DATA[9]~input_o ),
	.usb_DATA_10(\usb_DATA[10]~input_o ),
	.usb_DATA_11(\usb_DATA[11]~input_o ),
	.usb_DATA_12(\usb_DATA[12]~input_o ),
	.usb_DATA_13(\usb_DATA[13]~input_o ),
	.usb_DATA_14(\usb_DATA[14]~input_o ),
	.usb_DATA_15(\usb_DATA[15]~input_o ),
	.usb_INT(\usb_INT~input_o ));

usb_system_usb_system_all_switches all_switches(
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\all_switches|readdata[0]~q ),
	.readdata_1(\all_switches|readdata[1]~q ),
	.readdata_2(\all_switches|readdata[2]~q ),
	.readdata_3(\all_switches|readdata[3]~q ),
	.readdata_4(\all_switches|readdata[4]~q ),
	.readdata_5(\all_switches|readdata[5]~q ),
	.readdata_6(\all_switches|readdata[6]~q ),
	.readdata_7(\all_switches|readdata[7]~q ),
	.readdata_8(\all_switches|readdata[8]~q ),
	.readdata_9(\all_switches|readdata[9]~q ),
	.readdata_10(\all_switches|readdata[10]~q ),
	.readdata_11(\all_switches|readdata[11]~q ),
	.readdata_12(\all_switches|readdata[12]~q ),
	.readdata_13(\all_switches|readdata[13]~q ),
	.readdata_14(\all_switches|readdata[14]~q ),
	.readdata_15(\all_switches|readdata[15]~q ),
	.readdata_16(\all_switches|readdata[16]~q ),
	.readdata_17(\all_switches|readdata[17]~q ),
	.clk_clk(\clk_clk~input_o ),
	.all_switches_wire_export_0(\all_switches_wire_export[0]~input_o ),
	.all_switches_wire_export_1(\all_switches_wire_export[1]~input_o ),
	.all_switches_wire_export_2(\all_switches_wire_export[2]~input_o ),
	.all_switches_wire_export_3(\all_switches_wire_export[3]~input_o ),
	.all_switches_wire_export_4(\all_switches_wire_export[4]~input_o ),
	.all_switches_wire_export_5(\all_switches_wire_export[5]~input_o ),
	.all_switches_wire_export_6(\all_switches_wire_export[6]~input_o ),
	.all_switches_wire_export_7(\all_switches_wire_export[7]~input_o ),
	.all_switches_wire_export_8(\all_switches_wire_export[8]~input_o ),
	.all_switches_wire_export_9(\all_switches_wire_export[9]~input_o ),
	.all_switches_wire_export_10(\all_switches_wire_export[10]~input_o ),
	.all_switches_wire_export_11(\all_switches_wire_export[11]~input_o ),
	.all_switches_wire_export_12(\all_switches_wire_export[12]~input_o ),
	.all_switches_wire_export_13(\all_switches_wire_export[13]~input_o ),
	.all_switches_wire_export_14(\all_switches_wire_export[14]~input_o ),
	.all_switches_wire_export_15(\all_switches_wire_export[15]~input_o ),
	.all_switches_wire_export_16(\all_switches_wire_export[16]~input_o ),
	.all_switches_wire_export_17(\all_switches_wire_export[17]~input_o ));

usb_system_usb_system_jtag_uart jtag_uart(
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.tdo(\jtag_uart|usb_system_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller_002|r_sync_rst~q ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.sink_in_reset(\clock_crossing_io|cmd_fifo|sink_in_reset~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.uav_write(\mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest1(\jtag_uart|av_waitrequest~q ),
	.Equal9(\mm_interconnect_0|router|Equal9~1_combout ),
	.s0_cmd_valid(\clock_crossing_io|s0_cmd_valid~combout ),
	.sink_ready(\mm_interconnect_0|cmd_demux|sink_ready~11_combout ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.b_full(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.read_01(\jtag_uart|read_0~q ),
	.av_readdata_0(\jtag_uart|av_readdata[0]~1_combout ),
	.av_readdata_1(\jtag_uart|av_readdata[1]~2_combout ),
	.av_readdata_2(\jtag_uart|av_readdata[2]~3_combout ),
	.av_readdata_3(\jtag_uart|av_readdata[3]~4_combout ),
	.av_readdata_4(\jtag_uart|av_readdata[4]~5_combout ),
	.av_readdata_5(\jtag_uart|av_readdata[5]~6_combout ),
	.av_readdata_6(\jtag_uart|av_readdata[6]~7_combout ),
	.av_readdata_7(\jtag_uart|av_readdata[7]~8_combout ),
	.counter_reg_bit_3(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.b_full1(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_5(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.b_non_empty(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_31(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_21(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_01(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_11(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_41(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_51(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.ac1(\jtag_uart|ac~q ),
	.woverflow1(\jtag_uart|woverflow~q ),
	.rvalid1(\jtag_uart|rvalid~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

usb_system_usb_system_mm_interconnect_0 mm_interconnect_0(
	.wire_pll7_clk_0(\clocks|sd1|wire_pll7_clk[0] ),
	.W_alu_result_7(\cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_14(\cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_18(\cpu|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\cpu|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\cpu|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\cpu|cpu|W_alu_result[15]~q ),
	.W_alu_result_12(\cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_23(\cpu|cpu|W_alu_result[23]~q ),
	.W_alu_result_22(\cpu|cpu|W_alu_result[22]~q ),
	.W_alu_result_8(\cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_6(\cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_24(\cpu|cpu|W_alu_result[24]~q ),
	.W_alu_result_21(\cpu|cpu|W_alu_result[21]~q ),
	.W_alu_result_20(\cpu|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\cpu|cpu|W_alu_result[19]~q ),
	.W_alu_result_28(\cpu|cpu|W_alu_result[28]~q ),
	.W_alu_result_27(\cpu|cpu|W_alu_result[27]~q ),
	.W_alu_result_26(\cpu|cpu|W_alu_result[26]~q ),
	.W_alu_result_25(\cpu|cpu|W_alu_result[25]~q ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.readdata_0(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[0]~q ),
	.readdata_1(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_5(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_6(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[6]~q ),
	.d_writedata_24(\cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\cpu|cpu|d_writedata[26]~q ),
	.d_writedata_27(\cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\cpu|cpu|d_writedata[31]~q ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller_002|r_sync_rst~q ),
	.Equal3(\mm_interconnect_0|router|Equal3~4_combout ),
	.Equal6(\mm_interconnect_0|router|Equal6~0_combout ),
	.mem_used_1(\mm_interconnect_0|keycode_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\keycode|always0~0_combout ),
	.d_write(\cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|cpu_data_master_translator|write_accepted~q ),
	.wait_latency_counter_1(\mm_interconnect_0|keycode_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|keycode_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.mem_used_11(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always01(\led|always0~1_combout ),
	.wait_latency_counter_11(\mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ),
	.mem_used_12(\mm_interconnect_0|red_leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always02(\red_leds|always0~1_combout ),
	.wait_latency_counter_12(\mm_interconnect_0|red_leds_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_02(\mm_interconnect_0|red_leds_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_8(\cpu|cpu|d_writedata[8]~q ),
	.d_writedata_9(\cpu|cpu|d_writedata[9]~q ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.d_writedata_11(\cpu|cpu|d_writedata[11]~q ),
	.d_writedata_12(\cpu|cpu|d_writedata[12]~q ),
	.d_writedata_13(\cpu|cpu|d_writedata[13]~q ),
	.d_writedata_14(\cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\cpu|cpu|d_writedata[15]~q ),
	.d_writedata_16(\cpu|cpu|d_writedata[16]~q ),
	.d_writedata_17(\cpu|cpu|d_writedata[17]~q ),
	.entries_1(\sdram|the_usb_system_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_usb_system_sdram_input_efifo_module|entries[0]~q ),
	.altera_reset_synchronizer_int_chain_out1(\rst_controller_003|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.sink_in_reset(\clock_crossing_io|cmd_fifo|sink_in_reset~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|keycode_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|red_leds_s1_translator|read_latency_shift_reg[0]~q ),
	.out_valid(\clock_crossing_io|rsp_fifo|out_valid~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.read_latency_shift_reg_02(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\mm_interconnect_0|cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.read_latency_shift_reg_04(\mm_interconnect_0|led_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_05(\mm_interconnect_0|all_switches_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.mem_67_0(\mm_interconnect_0|sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_01(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_02(\mm_interconnect_0|clock_crossing_io_s0_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_03(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem[0][67]~q ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.mem_67_04(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_05(\mm_interconnect_0|keycode_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_06(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_07(\mm_interconnect_0|red_leds_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_08(\mm_interconnect_0|all_switches_s1_agent_rsp_fifo|mem[0][67]~q ),
	.out_valid1(\mm_interconnect_0|crosser_002|clock_xer|out_valid~combout ),
	.out_data_buffer_67(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[67]~q ),
	.av_ld_getting_data(\cpu|cpu|av_ld_getting_data~6_combout ),
	.waitrequest(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_13(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.uav_write(\mm_interconnect_0|cpu_data_master_translator|uav_write~0_combout ),
	.mem_used_14(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem_used[1]~q ),
	.full(\clock_crossing_io|cmd_fifo|full~q ),
	.F_pc_26(\cpu|cpu|F_pc[26]~q ),
	.F_pc_25(\cpu|cpu|F_pc[25]~q ),
	.F_pc_24(\cpu|cpu|F_pc[24]~q ),
	.F_pc_23(\cpu|cpu|F_pc[23]~q ),
	.F_pc_22(\cpu|cpu|F_pc[22]~q ),
	.F_pc_21(\cpu|cpu|F_pc[21]~q ),
	.F_pc_20(\cpu|cpu|F_pc[20]~q ),
	.F_pc_19(\cpu|cpu|F_pc[19]~q ),
	.F_pc_18(\cpu|cpu|F_pc[18]~q ),
	.F_pc_17(\cpu|cpu|F_pc[17]~q ),
	.F_pc_16(\cpu|cpu|F_pc[16]~q ),
	.F_pc_15(\cpu|cpu|F_pc[15]~q ),
	.F_pc_14(\cpu|cpu|F_pc[14]~q ),
	.F_pc_13(\cpu|cpu|F_pc[13]~q ),
	.F_pc_12(\cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\cpu|cpu|F_pc[11]~q ),
	.F_pc_10(\cpu|cpu|F_pc[10]~q ),
	.F_pc_9(\cpu|cpu|F_pc[9]~q ),
	.F_pc_8(\cpu|cpu|F_pc[8]~q ),
	.F_pc_7(\cpu|cpu|F_pc[7]~q ),
	.F_pc_5(\cpu|cpu|F_pc[5]~q ),
	.F_pc_6(\cpu|cpu|F_pc[6]~q ),
	.F_pc_4(\cpu|cpu|F_pc[4]~q ),
	.F_pc_1(\cpu|cpu|F_pc[1]~q ),
	.F_pc_3(\cpu|cpu|F_pc[3]~q ),
	.i_read(\cpu|cpu|i_read~q ),
	.F_pc_2(\cpu|cpu|F_pc[2]~q ),
	.mem_used_15(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\jtag_uart|av_waitrequest~q ),
	.Equal9(\mm_interconnect_0|router|Equal9~1_combout ),
	.cpu_data_master_waitrequest(\mm_interconnect_0|cpu_data_master_translator|av_waitrequest~1_combout ),
	.s0_cmd_valid(\clock_crossing_io|s0_cmd_valid~combout ),
	.WideOr11(\mm_interconnect_0|cmd_mux_003|WideOr1~combout ),
	.F_pc_0(\cpu|cpu|F_pc[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.mem(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem~0_combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.last_cycle(\mm_interconnect_0|cmd_mux_006|last_cycle~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.WideOr12(\mm_interconnect_0|cmd_mux_006|WideOr1~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_006|src_payload~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_006|src_data[68]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_006|src_data[48]~combout ),
	.src_data_62(\mm_interconnect_0|cmd_mux_006|src_data[62]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_006|src_data[49]~combout ),
	.src_data_51(\mm_interconnect_0|cmd_mux_006|src_data[51]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_006|src_data[50]~combout ),
	.src_data_53(\mm_interconnect_0|cmd_mux_006|src_data[53]~combout ),
	.src_data_52(\mm_interconnect_0|cmd_mux_006|src_data[52]~combout ),
	.src_data_55(\mm_interconnect_0|cmd_mux_006|src_data[55]~combout ),
	.src_data_54(\mm_interconnect_0|cmd_mux_006|src_data[54]~combout ),
	.src_data_57(\mm_interconnect_0|cmd_mux_006|src_data[57]~combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_006|src_data[56]~combout ),
	.src_data_59(\mm_interconnect_0|cmd_mux_006|src_data[59]~combout ),
	.src_data_58(\mm_interconnect_0|cmd_mux_006|src_data[58]~combout ),
	.src_data_61(\mm_interconnect_0|cmd_mux_006|src_data[61]~combout ),
	.src_data_60(\mm_interconnect_0|cmd_mux_006|src_data[60]~combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_006|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_006|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_006|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_006|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_006|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_006|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_006|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_006|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_006|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_006|src_data[47]~combout ),
	.out_data_buffer_32(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_321(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_33(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_331(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_34(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_341(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_35(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[35]~q ),
	.out_data_buffer_351(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[35]~q ),
	.sink_ready(\mm_interconnect_0|cmd_demux|sink_ready~11_combout ),
	.WideOr13(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.local_read(\mm_interconnect_0|cpu_debug_mem_slave_agent|local_read~0_combout ),
	.mem1(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem~1_combout ),
	.m0_write(\mm_interconnect_0|clock_crossing_io_s0_agent|m0_write~2_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.out_valid2(\mm_interconnect_0|crosser_003|clock_xer|out_valid~combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.WideOr14(\mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ),
	.av_readdatavalid(\mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~0_combout ),
	.av_readdatavalid1(\mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~1_combout ),
	.av_readdatavalid2(\mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~2_combout ),
	.hbreak_enabled(\cpu|cpu|hbreak_enabled~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[0]~q ),
	.av_readdata_pre_0(\mm_interconnect_0|clocks_pll_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|clocks_pll_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~2_combout ),
	.av_readdata_pre_3(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[4]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.out_payload_0(\clock_crossing_io|rsp_fifo|out_payload[0]~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.out_data_buffer_22(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[22]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.out_data_buffer_23(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_24(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.out_data_buffer_25(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_26(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.out_data_buffer_11(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[11]~q ),
	.av_readdata_pre_111(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_13(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[13]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~3_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[5]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_14(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_15(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[15]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_9(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[9]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_8(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[7]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[6]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_20(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.out_data_buffer_18(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.out_data_buffer_19(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[19]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.out_data_buffer_17(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[17]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~5_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.out_data_buffer_27(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_28(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.out_data_buffer_31(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_30(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.out_data_buffer_29(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[29]~q ),
	.mem2(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem~4_combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.out_payload_1(\clock_crossing_io|rsp_fifo|out_payload[1]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.out_payload_2(\clock_crossing_io|rsp_fifo|out_payload[2]~q ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~28_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~30_combout ),
	.out_payload_3(\clock_crossing_io|rsp_fifo|out_payload[3]~q ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[3]~34_combout ),
	.out_payload_4(\clock_crossing_io|rsp_fifo|out_payload[4]~q ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~37_combout ),
	.out_payload_5(\clock_crossing_io|rsp_fifo|out_payload[5]~q ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~41_combout ),
	.out_payload_6(\clock_crossing_io|rsp_fifo|out_payload[6]~q ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~45_combout ),
	.out_payload_7(\clock_crossing_io|rsp_fifo|out_payload[7]~q ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~49_combout ),
	.out_payload_8(\clock_crossing_io|rsp_fifo|out_payload[8]~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.readdata_01(\clocks|readdata[0]~1_combout ),
	.readdata_11(\clocks|readdata[1]~2_combout ),
	.readdata_4(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[4]~q ),
	.out_payload_9(\clock_crossing_io|rsp_fifo|out_payload[9]~q ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.out_payload_10(\clock_crossing_io|rsp_fifo|out_payload[10]~q ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~59_combout ),
	.out_payload_11(\clock_crossing_io|rsp_fifo|out_payload[11]~q ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.out_payload_12(\clock_crossing_io|rsp_fifo|out_payload[12]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~66_combout ),
	.out_payload_13(\clock_crossing_io|rsp_fifo|out_payload[13]~q ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~combout ),
	.out_payload_14(\clock_crossing_io|rsp_fifo|out_payload[14]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~72_combout ),
	.out_payload_15(\clock_crossing_io|rsp_fifo|out_payload[15]~q ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~78_combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~combout ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.d_byteenable_1(\cpu|cpu|d_byteenable[1]~q ),
	.d_byteenable_2(\cpu|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\cpu|cpu|d_byteenable[3]~q ),
	.b_full(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_payload8(\mm_interconnect_0|cmd_mux_006|src_payload~1_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_006|src_payload~2_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_006|src_payload~3_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_006|src_payload~4_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_006|src_payload~5_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_006|src_payload~6_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_006|src_payload~7_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_006|src_payload~8_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_006|src_payload~9_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_006|src_payload~10_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_006|src_payload~11_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_006|src_payload~12_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_006|src_payload~13_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_006|src_payload~14_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_006|src_payload~15_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_006|src_payload~16_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_006|src_payload~17_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_006|src_payload~18_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_006|src_payload~19_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_006|src_payload~20_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_006|src_payload~21_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_006|src_payload~22_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_006|src_payload~23_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_006|src_payload~24_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_006|src_payload~25_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_006|src_payload~26_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_006|src_payload~27_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_006|src_payload~28_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_006|src_payload~29_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_006|src_payload~30_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_006|src_payload~31_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_006|src_payload~32_combout ),
	.read_0(\jtag_uart|read_0~q ),
	.av_readdata_0(\jtag_uart|av_readdata[0]~1_combout ),
	.readdata_02(\led|readdata[0]~combout ),
	.readdata_03(\keycode|readdata[0]~combout ),
	.readdata_04(\all_switches|readdata[0]~q ),
	.readdata_05(\red_leds|readdata[0]~combout ),
	.readdata_22(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[22]~q ),
	.readdata_23(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[23]~q ),
	.readdata_24(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[26]~q ),
	.readdata_111(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[11]~q ),
	.readdata_13(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[13]~q ),
	.readdata_16(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_12(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[12]~q ),
	.readdata_14(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[14]~q ),
	.readdata_15(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[15]~q ),
	.readdata_10(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[10]~q ),
	.readdata_9(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[9]~q ),
	.readdata_8(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[8]~q ),
	.readdata_7(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_20(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[20]~q ),
	.readdata_18(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[18]~q ),
	.readdata_19(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[19]~q ),
	.readdata_17(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[17]~q ),
	.src_payload40(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.readdata_21(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[21]~q ),
	.src_payload41(\mm_interconnect_0|rsp_mux|src_payload~12_combout ),
	.readdata_27(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[27]~q ),
	.src_payload42(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.src_payload43(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.src_payload44(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.src_payload45(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.out_data_buffer_241(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[24]~q ),
	.readdata_28(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[28]~q ),
	.out_data_buffer_281(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_271(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[27]~q ),
	.readdata_31(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[31]~q ),
	.out_data_buffer_261(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[26]~q ),
	.readdata_30(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[30]~q ),
	.out_data_buffer_251(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[25]~q ),
	.readdata_29(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[29]~q ),
	.av_readdata_1(\jtag_uart|av_readdata[1]~2_combout ),
	.readdata_110(\led|readdata[1]~combout ),
	.readdata_112(\keycode|readdata[1]~combout ),
	.readdata_113(\all_switches|readdata[1]~q ),
	.readdata_114(\red_leds|readdata[1]~combout ),
	.av_readdata_2(\jtag_uart|av_readdata[2]~3_combout ),
	.readdata_210(\led|readdata[2]~combout ),
	.readdata_211(\keycode|readdata[2]~combout ),
	.readdata_212(\all_switches|readdata[2]~q ),
	.readdata_213(\red_leds|readdata[2]~combout ),
	.readdata_32(\all_switches|readdata[3]~q ),
	.readdata_33(\red_leds|readdata[3]~combout ),
	.av_readdata_3(\jtag_uart|av_readdata[3]~4_combout ),
	.readdata_34(\led|readdata[3]~combout ),
	.readdata_35(\keycode|readdata[3]~combout ),
	.av_readdata_4(\jtag_uart|av_readdata[4]~5_combout ),
	.readdata_41(\led|readdata[4]~combout ),
	.readdata_42(\keycode|readdata[4]~combout ),
	.readdata_43(\all_switches|readdata[4]~q ),
	.readdata_44(\red_leds|readdata[4]~combout ),
	.av_readdata_5(\jtag_uart|av_readdata[5]~6_combout ),
	.readdata_51(\led|readdata[5]~combout ),
	.readdata_52(\keycode|readdata[5]~combout ),
	.readdata_53(\all_switches|readdata[5]~q ),
	.readdata_54(\red_leds|readdata[5]~combout ),
	.av_readdata_6(\jtag_uart|av_readdata[6]~7_combout ),
	.readdata_61(\led|readdata[6]~combout ),
	.readdata_62(\keycode|readdata[6]~combout ),
	.readdata_63(\all_switches|readdata[6]~q ),
	.readdata_64(\red_leds|readdata[6]~combout ),
	.av_readdata_7(\jtag_uart|av_readdata[7]~8_combout ),
	.readdata_71(\led|readdata[7]~combout ),
	.readdata_72(\keycode|readdata[7]~combout ),
	.readdata_73(\all_switches|readdata[7]~q ),
	.readdata_74(\red_leds|readdata[7]~combout ),
	.readdata_81(\all_switches|readdata[8]~q ),
	.readdata_82(\red_leds|readdata[8]~combout ),
	.counter_reg_bit_3(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.b_full1(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_5(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart|the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.b_non_empty(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_31(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_21(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_01(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_11(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_41(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_51(\jtag_uart|the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.readdata_91(\all_switches|readdata[9]~q ),
	.readdata_92(\red_leds|readdata[9]~combout ),
	.ac(\jtag_uart|ac~q ),
	.readdata_101(\all_switches|readdata[10]~q ),
	.readdata_102(\red_leds|readdata[10]~combout ),
	.readdata_115(\all_switches|readdata[11]~q ),
	.readdata_116(\red_leds|readdata[11]~combout ),
	.readdata_121(\all_switches|readdata[12]~q ),
	.readdata_122(\red_leds|readdata[12]~combout ),
	.readdata_131(\all_switches|readdata[13]~q ),
	.readdata_132(\red_leds|readdata[13]~combout ),
	.woverflow(\jtag_uart|woverflow~q ),
	.readdata_141(\all_switches|readdata[14]~q ),
	.readdata_142(\red_leds|readdata[14]~combout ),
	.readdata_151(\all_switches|readdata[15]~q ),
	.readdata_152(\red_leds|readdata[15]~combout ),
	.rvalid(\jtag_uart|rvalid~q ),
	.readdata_161(\all_switches|readdata[16]~q ),
	.readdata_162(\red_leds|readdata[16]~combout ),
	.readdata_171(\all_switches|readdata[17]~q ),
	.readdata_172(\red_leds|readdata[17]~combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_382(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_392(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.out_data_buffer_311(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_301(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_291(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[29]~q ),
	.src_payload48(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.za_valid(\sdram|za_valid~q ),
	.src_payload51(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.d_writedata_18(\cpu|cpu|d_writedata[18]~q ),
	.d_writedata_19(\cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\cpu|cpu|d_writedata[20]~q ),
	.d_writedata_21(\cpu|cpu|d_writedata[21]~q ),
	.d_writedata_22(\cpu|cpu|d_writedata[22]~q ),
	.d_writedata_23(\cpu|cpu|d_writedata[23]~q ),
	.src_payload52(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload56(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload62(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload65(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload66(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload67(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload74(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload75(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload76(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload77(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.za_data_0(\sdram|za_data[0]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.za_data_22(\sdram|za_data[22]~q ),
	.za_data_23(\sdram|za_data[23]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.za_data_16(\sdram|za_data[16]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.za_data_20(\sdram|za_data[20]~q ),
	.za_data_18(\sdram|za_data[18]~q ),
	.za_data_19(\sdram|za_data[19]~q ),
	.za_data_17(\sdram|za_data[17]~q ),
	.za_data_21(\sdram|za_data[21]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.m0_write1(\mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ),
	.m0_read(\mm_interconnect_0|clock_crossing_io_s0_agent|m0_read~2_combout ),
	.m0_write2(\mm_interconnect_0|clock_crossing_io_s0_agent|m0_write~3_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~84_combout ),
	.src_data_410(\mm_interconnect_0|rsp_mux|src_data[4]~85_combout ),
	.src_data_510(\mm_interconnect_0|rsp_mux|src_data[5]~86_combout ),
	.src_data_63(\mm_interconnect_0|rsp_mux|src_data[6]~87_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux|src_data[7]~88_combout ),
	.clk_clk(\clk_clk~input_o ));

usb_system_usb_system_sdram sdram(
	.wire_pll7_clk_0(\clocks|sd1|wire_pll7_clk[0] ),
	.m_addr_0(\sdram|m_addr[0]~q ),
	.m_addr_1(\sdram|m_addr[1]~q ),
	.m_addr_2(\sdram|m_addr[2]~q ),
	.m_addr_3(\sdram|m_addr[3]~q ),
	.m_addr_4(\sdram|m_addr[4]~q ),
	.m_addr_5(\sdram|m_addr[5]~q ),
	.m_addr_6(\sdram|m_addr[6]~q ),
	.m_addr_7(\sdram|m_addr[7]~q ),
	.m_addr_8(\sdram|m_addr[8]~q ),
	.m_addr_9(\sdram|m_addr[9]~q ),
	.oe1(\sdram|oe~q ),
	.m_addr_10(\sdram|m_addr[10]~q ),
	.m_addr_11(\sdram|m_addr[11]~q ),
	.m_addr_12(\sdram|m_addr[12]~q ),
	.m_bank_0(\sdram|m_bank[0]~q ),
	.m_bank_1(\sdram|m_bank[1]~q ),
	.m_cmd_1(\sdram|m_cmd[1]~q ),
	.m_cmd_3(\sdram|m_cmd[3]~q ),
	.m_dqm_0(\sdram|m_dqm[0]~q ),
	.m_dqm_1(\sdram|m_dqm[1]~q ),
	.m_dqm_2(\sdram|m_dqm[2]~q ),
	.m_dqm_3(\sdram|m_dqm[3]~q ),
	.m_cmd_2(\sdram|m_cmd[2]~q ),
	.m_cmd_0(\sdram|m_cmd[0]~q ),
	.entries_1(\sdram|the_usb_system_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_usb_system_sdram_input_efifo_module|entries[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_003|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.last_cycle(\mm_interconnect_0|cmd_mux_006|last_cycle~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_006|WideOr1~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_006|src_payload~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_006|src_data[68]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_006|src_data[48]~combout ),
	.src_data_62(\mm_interconnect_0|cmd_mux_006|src_data[62]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_006|src_data[49]~combout ),
	.src_data_51(\mm_interconnect_0|cmd_mux_006|src_data[51]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_006|src_data[50]~combout ),
	.src_data_53(\mm_interconnect_0|cmd_mux_006|src_data[53]~combout ),
	.src_data_52(\mm_interconnect_0|cmd_mux_006|src_data[52]~combout ),
	.src_data_55(\mm_interconnect_0|cmd_mux_006|src_data[55]~combout ),
	.src_data_54(\mm_interconnect_0|cmd_mux_006|src_data[54]~combout ),
	.src_data_57(\mm_interconnect_0|cmd_mux_006|src_data[57]~combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_006|src_data[56]~combout ),
	.src_data_59(\mm_interconnect_0|cmd_mux_006|src_data[59]~combout ),
	.src_data_58(\mm_interconnect_0|cmd_mux_006|src_data[58]~combout ),
	.src_data_61(\mm_interconnect_0|cmd_mux_006|src_data[61]~combout ),
	.src_data_60(\mm_interconnect_0|cmd_mux_006|src_data[60]~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_006|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_006|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_006|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_006|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_006|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_006|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_006|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_006|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_006|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_006|src_data[47]~combout ),
	.out_data_buffer_32(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_321(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_33(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_331(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_34(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_341(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_35(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[35]~q ),
	.out_data_buffer_351(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[35]~q ),
	.m_data_0(\sdram|m_data[0]~q ),
	.m_data_1(\sdram|m_data[1]~q ),
	.m_data_2(\sdram|m_data[2]~q ),
	.m_data_3(\sdram|m_data[3]~q ),
	.m_data_4(\sdram|m_data[4]~q ),
	.m_data_5(\sdram|m_data[5]~q ),
	.m_data_6(\sdram|m_data[6]~q ),
	.m_data_7(\sdram|m_data[7]~q ),
	.m_data_8(\sdram|m_data[8]~q ),
	.m_data_9(\sdram|m_data[9]~q ),
	.m_data_10(\sdram|m_data[10]~q ),
	.m_data_11(\sdram|m_data[11]~q ),
	.m_data_12(\sdram|m_data[12]~q ),
	.m_data_13(\sdram|m_data[13]~q ),
	.m_data_14(\sdram|m_data[14]~q ),
	.m_data_15(\sdram|m_data[15]~q ),
	.m_data_16(\sdram|m_data[16]~q ),
	.m_data_17(\sdram|m_data[17]~q ),
	.m_data_18(\sdram|m_data[18]~q ),
	.m_data_19(\sdram|m_data[19]~q ),
	.m_data_20(\sdram|m_data[20]~q ),
	.m_data_21(\sdram|m_data[21]~q ),
	.m_data_22(\sdram|m_data[22]~q ),
	.m_data_23(\sdram|m_data[23]~q ),
	.m_data_24(\sdram|m_data[24]~q ),
	.m_data_25(\sdram|m_data[25]~q ),
	.m_data_26(\sdram|m_data[26]~q ),
	.m_data_27(\sdram|m_data[27]~q ),
	.m_data_28(\sdram|m_data[28]~q ),
	.m_data_29(\sdram|m_data[29]~q ),
	.m_data_30(\sdram|m_data[30]~q ),
	.m_data_31(\sdram|m_data[31]~q ),
	.src_payload1(\mm_interconnect_0|cmd_mux_006|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_006|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_006|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_006|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_006|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_006|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_006|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_006|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_006|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_006|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_006|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_006|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_006|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_006|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_006|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_006|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_006|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_006|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_006|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_006|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_006|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_006|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_006|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_006|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_006|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_006|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_006|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_006|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_006|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_006|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_006|src_payload~31_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_006|src_payload~32_combout ),
	.za_valid1(\sdram|za_valid~q ),
	.za_data_0(\sdram|za_data[0]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.za_data_22(\sdram|za_data[22]~q ),
	.za_data_23(\sdram|za_data[23]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.za_data_16(\sdram|za_data[16]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.za_data_20(\sdram|za_data[20]~q ),
	.za_data_18(\sdram|za_data[18]~q ),
	.za_data_19(\sdram|za_data[19]~q ),
	.za_data_17(\sdram|za_data[17]~q ),
	.za_data_21(\sdram|za_data[21]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.m0_write(\mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ),
	.sdram_wire_dq_0(\sdram_wire_dq[0]~input_o ),
	.sdram_wire_dq_1(\sdram_wire_dq[1]~input_o ),
	.sdram_wire_dq_2(\sdram_wire_dq[2]~input_o ),
	.sdram_wire_dq_3(\sdram_wire_dq[3]~input_o ),
	.sdram_wire_dq_4(\sdram_wire_dq[4]~input_o ),
	.sdram_wire_dq_5(\sdram_wire_dq[5]~input_o ),
	.sdram_wire_dq_6(\sdram_wire_dq[6]~input_o ),
	.sdram_wire_dq_7(\sdram_wire_dq[7]~input_o ),
	.sdram_wire_dq_8(\sdram_wire_dq[8]~input_o ),
	.sdram_wire_dq_9(\sdram_wire_dq[9]~input_o ),
	.sdram_wire_dq_10(\sdram_wire_dq[10]~input_o ),
	.sdram_wire_dq_11(\sdram_wire_dq[11]~input_o ),
	.sdram_wire_dq_12(\sdram_wire_dq[12]~input_o ),
	.sdram_wire_dq_13(\sdram_wire_dq[13]~input_o ),
	.sdram_wire_dq_14(\sdram_wire_dq[14]~input_o ),
	.sdram_wire_dq_15(\sdram_wire_dq[15]~input_o ),
	.sdram_wire_dq_16(\sdram_wire_dq[16]~input_o ),
	.sdram_wire_dq_17(\sdram_wire_dq[17]~input_o ),
	.sdram_wire_dq_18(\sdram_wire_dq[18]~input_o ),
	.sdram_wire_dq_19(\sdram_wire_dq[19]~input_o ),
	.sdram_wire_dq_20(\sdram_wire_dq[20]~input_o ),
	.sdram_wire_dq_21(\sdram_wire_dq[21]~input_o ),
	.sdram_wire_dq_22(\sdram_wire_dq[22]~input_o ),
	.sdram_wire_dq_23(\sdram_wire_dq[23]~input_o ),
	.sdram_wire_dq_24(\sdram_wire_dq[24]~input_o ),
	.sdram_wire_dq_25(\sdram_wire_dq[25]~input_o ),
	.sdram_wire_dq_26(\sdram_wire_dq[26]~input_o ),
	.sdram_wire_dq_27(\sdram_wire_dq[27]~input_o ),
	.sdram_wire_dq_28(\sdram_wire_dq[28]~input_o ),
	.sdram_wire_dq_29(\sdram_wire_dq[29]~input_o ),
	.sdram_wire_dq_30(\sdram_wire_dq[30]~input_o ),
	.sdram_wire_dq_31(\sdram_wire_dq[31]~input_o ));

usb_system_usb_system_red_leds red_leds(
	.W_alu_result_7(\cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.data_out_0(\red_leds|data_out[0]~q ),
	.data_out_1(\red_leds|data_out[1]~q ),
	.data_out_2(\red_leds|data_out[2]~q ),
	.data_out_3(\red_leds|data_out[3]~q ),
	.data_out_4(\red_leds|data_out[4]~q ),
	.data_out_5(\red_leds|data_out[5]~q ),
	.data_out_6(\red_leds|data_out[6]~q ),
	.data_out_7(\red_leds|data_out[7]~q ),
	.data_out_8(\red_leds|data_out[8]~q ),
	.data_out_9(\red_leds|data_out[9]~q ),
	.data_out_10(\red_leds|data_out[10]~q ),
	.data_out_11(\red_leds|data_out[11]~q ),
	.data_out_12(\red_leds|data_out[12]~q ),
	.data_out_13(\red_leds|data_out[13]~q ),
	.data_out_14(\red_leds|data_out[14]~q ),
	.data_out_15(\red_leds|data_out[15]~q ),
	.data_out_16(\red_leds|data_out[16]~q ),
	.data_out_17(\red_leds|data_out[17]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|cpu|d_writedata[17]~q ,\cpu|cpu|d_writedata[16]~q ,\cpu|cpu|d_writedata[15]~q ,\cpu|cpu|d_writedata[14]~q ,\cpu|cpu|d_writedata[13]~q ,\cpu|cpu|d_writedata[12]~q ,\cpu|cpu|d_writedata[11]~q ,
\cpu|cpu|d_writedata[10]~q ,\cpu|cpu|d_writedata[9]~q ,\cpu|cpu|d_writedata[8]~q ,\cpu|cpu|d_writedata[7]~q ,\cpu|cpu|d_writedata[6]~q ,\cpu|cpu|d_writedata[5]~q ,\cpu|cpu|d_writedata[4]~q ,\cpu|cpu|d_writedata[3]~q ,\cpu|cpu|d_writedata[2]~q ,
\cpu|cpu|d_writedata[1]~q ,\cpu|cpu|d_writedata[0]~q }),
	.Equal3(\mm_interconnect_0|router|Equal3~4_combout ),
	.always0(\keycode|always0~1_combout ),
	.reset_n(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.mem_used_1(\mm_interconnect_0|red_leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always01(\red_leds|always0~1_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|red_leds_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|red_leds_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\red_leds|readdata[0]~combout ),
	.readdata_1(\red_leds|readdata[1]~combout ),
	.readdata_2(\red_leds|readdata[2]~combout ),
	.readdata_3(\red_leds|readdata[3]~combout ),
	.readdata_4(\red_leds|readdata[4]~combout ),
	.readdata_5(\red_leds|readdata[5]~combout ),
	.readdata_6(\red_leds|readdata[6]~combout ),
	.readdata_7(\red_leds|readdata[7]~combout ),
	.readdata_8(\red_leds|readdata[8]~combout ),
	.readdata_9(\red_leds|readdata[9]~combout ),
	.readdata_10(\red_leds|readdata[10]~combout ),
	.readdata_11(\red_leds|readdata[11]~combout ),
	.readdata_12(\red_leds|readdata[12]~combout ),
	.readdata_13(\red_leds|readdata[13]~combout ),
	.readdata_14(\red_leds|readdata[14]~combout ),
	.readdata_15(\red_leds|readdata[15]~combout ),
	.readdata_16(\red_leds|readdata[16]~combout ),
	.readdata_17(\red_leds|readdata[17]~combout ),
	.clk(\clk_clk~input_o ));

usb_system_usb_system_keycode_1 led(
	.W_alu_result_7(\cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.data_out_0(\led|data_out[0]~q ),
	.data_out_1(\led|data_out[1]~q ),
	.data_out_2(\led|data_out[2]~q ),
	.data_out_3(\led|data_out[3]~q ),
	.data_out_4(\led|data_out[4]~q ),
	.data_out_5(\led|data_out[5]~q ),
	.data_out_6(\led|data_out[6]~q ),
	.data_out_7(\led|data_out[7]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|cpu|d_writedata[7]~q ,\cpu|cpu|d_writedata[6]~q ,\cpu|cpu|d_writedata[5]~q ,\cpu|cpu|d_writedata[4]~q ,\cpu|cpu|d_writedata[3]~q ,\cpu|cpu|d_writedata[2]~q ,\cpu|cpu|d_writedata[1]~q ,
\cpu|cpu|d_writedata[0]~q }),
	.Equal3(\mm_interconnect_0|router|Equal3~4_combout ),
	.always0(\keycode|always0~1_combout ),
	.reset_n(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.mem_used_1(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always01(\led|always0~1_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|led_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|led_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\led|readdata[0]~combout ),
	.readdata_1(\led|readdata[1]~combout ),
	.readdata_2(\led|readdata[2]~combout ),
	.readdata_3(\led|readdata[3]~combout ),
	.readdata_4(\led|readdata[4]~combout ),
	.readdata_5(\led|readdata[5]~combout ),
	.readdata_6(\led|readdata[6]~combout ),
	.readdata_7(\led|readdata[7]~combout ),
	.clk(\clk_clk~input_o ));

usb_system_usb_system_keycode keycode(
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.data_out_0(\keycode|data_out[0]~q ),
	.data_out_1(\keycode|data_out[1]~q ),
	.data_out_2(\keycode|data_out[2]~q ),
	.data_out_3(\keycode|data_out[3]~q ),
	.data_out_4(\keycode|data_out[4]~q ),
	.data_out_5(\keycode|data_out[5]~q ),
	.data_out_6(\keycode|data_out[6]~q ),
	.data_out_7(\keycode|data_out[7]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|cpu|d_writedata[7]~q ,\cpu|cpu|d_writedata[6]~q ,\cpu|cpu|d_writedata[5]~q ,\cpu|cpu|d_writedata[4]~q ,\cpu|cpu|d_writedata[3]~q ,\cpu|cpu|d_writedata[2]~q ,\cpu|cpu|d_writedata[1]~q ,
\cpu|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller_002|r_sync_rst~q ),
	.Equal6(\mm_interconnect_0|router|Equal6~0_combout ),
	.mem_used_1(\mm_interconnect_0|keycode_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\keycode|always0~0_combout ),
	.d_write(\cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|cpu_data_master_translator|write_accepted~q ),
	.always01(\keycode|always0~1_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|keycode_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|keycode_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\keycode|readdata[0]~combout ),
	.readdata_1(\keycode|readdata[1]~combout ),
	.readdata_2(\keycode|readdata[2]~combout ),
	.readdata_3(\keycode|readdata[3]~combout ),
	.readdata_4(\keycode|readdata[4]~combout ),
	.readdata_5(\keycode|readdata[5]~combout ),
	.readdata_6(\keycode|readdata[6]~combout ),
	.readdata_7(\keycode|readdata[7]~combout ),
	.clk(\clk_clk~input_o ));

usb_system_usb_system_cpu cpu(
	.sr_0(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.W_alu_result_7(\cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_14(\cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_18(\cpu|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\cpu|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\cpu|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\cpu|cpu|W_alu_result[15]~q ),
	.W_alu_result_12(\cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_11(\cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_23(\cpu|cpu|W_alu_result[23]~q ),
	.W_alu_result_22(\cpu|cpu|W_alu_result[22]~q ),
	.W_alu_result_8(\cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_6(\cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_24(\cpu|cpu|W_alu_result[24]~q ),
	.W_alu_result_21(\cpu|cpu|W_alu_result[21]~q ),
	.W_alu_result_20(\cpu|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\cpu|cpu|W_alu_result[19]~q ),
	.W_alu_result_28(\cpu|cpu|W_alu_result[28]~q ),
	.W_alu_result_27(\cpu|cpu|W_alu_result[27]~q ),
	.W_alu_result_26(\cpu|cpu|W_alu_result[26]~q ),
	.W_alu_result_25(\cpu|cpu|W_alu_result[25]~q ),
	.W_alu_result_4(\cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_5(\cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.readdata_0(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[0]~q ),
	.readdata_1(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_5(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_6(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[6]~q ),
	.d_writedata_24(\cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\cpu|cpu|d_writedata[26]~q ),
	.d_writedata_27(\cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\cpu|cpu|d_writedata[31]~q ),
	.ir_out_0(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller_002|r_sync_rst~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.d_writedata_8(\cpu|cpu|d_writedata[8]~q ),
	.d_writedata_9(\cpu|cpu|d_writedata[9]~q ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.d_writedata_11(\cpu|cpu|d_writedata[11]~q ),
	.d_writedata_12(\cpu|cpu|d_writedata[12]~q ),
	.d_writedata_13(\cpu|cpu|d_writedata[13]~q ),
	.d_writedata_14(\cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\cpu|cpu|d_writedata[15]~q ),
	.d_writedata_16(\cpu|cpu|d_writedata[16]~q ),
	.d_writedata_17(\cpu|cpu|d_writedata[17]~q ),
	.debug_reset_request(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_oci_debug|resetrequest~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|keycode_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|red_leds_s1_translator|read_latency_shift_reg[0]~q ),
	.out_valid(\clock_crossing_io|rsp_fifo|out_valid~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.read_latency_shift_reg_02(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\mm_interconnect_0|cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.read_latency_shift_reg_04(\mm_interconnect_0|led_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_05(\mm_interconnect_0|all_switches_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.mem_67_0(\mm_interconnect_0|sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_01(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_02(\mm_interconnect_0|clock_crossing_io_s0_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_03(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem[0][67]~q ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.mem_67_04(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_05(\mm_interconnect_0|keycode_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_06(\mm_interconnect_0|led_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_07(\mm_interconnect_0|red_leds_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_08(\mm_interconnect_0|all_switches_s1_agent_rsp_fifo|mem[0][67]~q ),
	.out_valid1(\mm_interconnect_0|crosser_002|clock_xer|out_valid~combout ),
	.out_data_buffer_67(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[67]~q ),
	.av_ld_getting_data(\cpu|cpu|av_ld_getting_data~6_combout ),
	.debug_mem_slave_waitrequest(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.F_pc_26(\cpu|cpu|F_pc[26]~q ),
	.F_pc_25(\cpu|cpu|F_pc[25]~q ),
	.F_pc_24(\cpu|cpu|F_pc[24]~q ),
	.F_pc_23(\cpu|cpu|F_pc[23]~q ),
	.F_pc_22(\cpu|cpu|F_pc[22]~q ),
	.F_pc_21(\cpu|cpu|F_pc[21]~q ),
	.F_pc_20(\cpu|cpu|F_pc[20]~q ),
	.F_pc_19(\cpu|cpu|F_pc[19]~q ),
	.F_pc_18(\cpu|cpu|F_pc[18]~q ),
	.F_pc_17(\cpu|cpu|F_pc[17]~q ),
	.F_pc_16(\cpu|cpu|F_pc[16]~q ),
	.F_pc_15(\cpu|cpu|F_pc[15]~q ),
	.F_pc_14(\cpu|cpu|F_pc[14]~q ),
	.F_pc_13(\cpu|cpu|F_pc[13]~q ),
	.F_pc_12(\cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\cpu|cpu|F_pc[11]~q ),
	.F_pc_10(\cpu|cpu|F_pc[10]~q ),
	.F_pc_9(\cpu|cpu|F_pc[9]~q ),
	.F_pc_8(\cpu|cpu|F_pc[8]~q ),
	.F_pc_7(\cpu|cpu|F_pc[7]~q ),
	.F_pc_5(\cpu|cpu|F_pc[5]~q ),
	.F_pc_6(\cpu|cpu|F_pc[6]~q ),
	.F_pc_4(\cpu|cpu|F_pc[4]~q ),
	.F_pc_1(\cpu|cpu|F_pc[1]~q ),
	.F_pc_3(\cpu|cpu|F_pc[3]~q ),
	.i_read(\cpu|cpu|i_read~q ),
	.F_pc_2(\cpu|cpu|F_pc[2]~q ),
	.av_waitrequest(\mm_interconnect_0|cpu_data_master_translator|av_waitrequest~1_combout ),
	.F_pc_0(\cpu|cpu|F_pc[0]~q ),
	.WideOr11(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.local_read(\mm_interconnect_0|cpu_debug_mem_slave_agent|local_read~0_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.out_valid2(\mm_interconnect_0|crosser_003|clock_xer|out_valid~combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.WideOr12(\mm_interconnect_0|rsp_mux_001|WideOr1~0_combout ),
	.av_readdatavalid(\mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~0_combout ),
	.av_readdatavalid1(\mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~1_combout ),
	.av_readdatavalid2(\mm_interconnect_0|cpu_instruction_master_agent|av_readdatavalid~2_combout ),
	.hbreak_enabled(\cpu|cpu|hbreak_enabled~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[0]~q ),
	.av_readdata_pre_0(\mm_interconnect_0|clocks_pll_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|clocks_pll_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~2_combout ),
	.av_readdata_pre_3(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[4]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.out_data_buffer_22(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[22]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.out_data_buffer_23(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_24(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.out_data_buffer_25(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_26(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.out_data_buffer_11(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[11]~q ),
	.av_readdata_pre_111(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_13(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[13]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~3_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[5]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_14(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_15(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[15]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_9(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[9]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_8(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[7]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[6]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_20(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.out_data_buffer_18(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.out_data_buffer_19(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[19]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.out_data_buffer_17(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[17]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~5_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.out_data_buffer_27(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_28(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.out_data_buffer_31(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_30(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.out_data_buffer_29(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[29]~q ),
	.mem(\mm_interconnect_0|cpu_debug_mem_slave_agent_rsp_fifo|mem~4_combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~28_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~30_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[3]~34_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~37_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~41_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~45_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~49_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.dreg_1(\irq_synchronizer|sync|sync[0].u|dreg[1]~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.readdata_4(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[4]~q ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~59_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~66_combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~72_combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~78_combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~combout ),
	.d_byteenable_0(\cpu|cpu|d_byteenable[0]~q ),
	.d_byteenable_1(\cpu|cpu|d_byteenable[1]~q ),
	.d_byteenable_2(\cpu|cpu|d_byteenable[2]~q ),
	.d_byteenable_3(\cpu|cpu|d_byteenable[3]~q ),
	.r_early_rst(\rst_controller_002|r_early_rst~q ),
	.readdata_22(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[22]~q ),
	.readdata_23(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[23]~q ),
	.readdata_24(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[26]~q ),
	.readdata_11(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[11]~q ),
	.readdata_13(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[13]~q ),
	.readdata_16(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_12(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[12]~q ),
	.readdata_14(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[14]~q ),
	.readdata_15(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[15]~q ),
	.readdata_10(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[10]~q ),
	.readdata_9(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[9]~q ),
	.readdata_8(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[8]~q ),
	.readdata_7(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_20(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[20]~q ),
	.readdata_18(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[18]~q ),
	.readdata_19(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[19]~q ),
	.readdata_17(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[17]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.readdata_21(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[21]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~12_combout ),
	.readdata_27(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[27]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.out_data_buffer_241(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[24]~q ),
	.readdata_28(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[28]~q ),
	.out_data_buffer_281(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_271(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[27]~q ),
	.readdata_31(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[31]~q ),
	.out_data_buffer_261(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[26]~q ),
	.readdata_30(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[30]~q ),
	.out_data_buffer_251(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[25]~q ),
	.readdata_29(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|readdata[29]~q ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.out_data_buffer_311(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_301(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_291(\mm_interconnect_0|crosser_002|clock_xer|out_data_buffer[29]~q ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.d_writedata_18(\cpu|cpu|d_writedata[18]~q ),
	.d_writedata_19(\cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\cpu|cpu|d_writedata[20]~q ),
	.d_writedata_21(\cpu|cpu|d_writedata[21]~q ),
	.d_writedata_22(\cpu|cpu|d_writedata[22]~q ),
	.d_writedata_23(\cpu|cpu|d_writedata[23]~q ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~84_combout ),
	.src_data_47(\mm_interconnect_0|rsp_mux|src_data[4]~85_combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux|src_data[5]~86_combout ),
	.src_data_61(\mm_interconnect_0|rsp_mux|src_data[6]~87_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux|src_data[7]~88_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

usb_system_usb_system_clocks clocks(
	.wire_pll7_clk_0(\clocks|sd1|wire_pll7_clk[0] ),
	.wire_pll7_clk_1(\clocks|sd1|wire_pll7_clk[1] ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.reset(\rst_controller_002|r_sync_rst~q ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.mem_used_1(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_003|WideOr1~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.mem(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem~0_combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.mem1(\mm_interconnect_0|clocks_pll_slave_agent_rsp_fifo|mem~1_combout ),
	.readdata_0(\clocks|readdata[0]~1_combout ),
	.readdata_1(\clocks|readdata[1]~2_combout ),
	.clk_clk(\clk_clk~input_o ));

usb_system_altera_avalon_mm_clock_crossing_bridge clock_crossing_io(
	.wire_pll7_clk_1(\clocks|sd1|wire_pll7_clk[1] ),
	.W_alu_result_2(\cpu|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\cpu|cpu|W_alu_result[3]~q ),
	.m0_reset(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.d_writedata_0(\cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller_002|r_sync_rst~q ),
	.d_write(\cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|cpu_data_master_translator|write_accepted~q ),
	.d_writedata_1(\cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\cpu|cpu|d_writedata[7]~q ),
	.d_writedata_8(\cpu|cpu|d_writedata[8]~q ),
	.d_writedata_9(\cpu|cpu|d_writedata[9]~q ),
	.d_writedata_10(\cpu|cpu|d_writedata[10]~q ),
	.d_writedata_11(\cpu|cpu|d_writedata[11]~q ),
	.d_writedata_12(\cpu|cpu|d_writedata[12]~q ),
	.d_writedata_13(\cpu|cpu|d_writedata[13]~q ),
	.d_writedata_14(\cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\cpu|cpu|d_writedata[15]~q ),
	.out_payload_42(\clock_crossing_io|cmd_fifo|out_payload[42]~q ),
	.out_payload_43(\clock_crossing_io|cmd_fifo|out_payload[43]~q ),
	.out_valid(\clock_crossing_io|cmd_fifo|out_valid~q ),
	.m0_read(\clock_crossing_io|m0_read~0_combout ),
	.out_payload_37(\clock_crossing_io|cmd_fifo|out_payload[37]~q ),
	.sink_in_reset(\clock_crossing_io|cmd_fifo|sink_in_reset~q ),
	.d_read(\cpu|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.out_valid1(\clock_crossing_io|rsp_fifo|out_valid~q ),
	.full(\clock_crossing_io|cmd_fifo|full~q ),
	.s0_cmd_valid1(\clock_crossing_io|s0_cmd_valid~combout ),
	.waitrequest_reset_override(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|waitrequest_reset_override~q ),
	.av_waitrequest_generated(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_waitrequest_generated~1_combout ),
	.m0_write(\mm_interconnect_0|clock_crossing_io_s0_agent|m0_write~2_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|read_latency_shift_reg[0]~q ),
	.out_payload_5(\clock_crossing_io|cmd_fifo|out_payload[5]~q ),
	.out_payload_6(\clock_crossing_io|cmd_fifo|out_payload[6]~q ),
	.out_payload_7(\clock_crossing_io|cmd_fifo|out_payload[7]~q ),
	.out_payload_8(\clock_crossing_io|cmd_fifo|out_payload[8]~q ),
	.out_payload_9(\clock_crossing_io|cmd_fifo|out_payload[9]~q ),
	.out_payload_10(\clock_crossing_io|cmd_fifo|out_payload[10]~q ),
	.out_payload_11(\clock_crossing_io|cmd_fifo|out_payload[11]~q ),
	.out_payload_12(\clock_crossing_io|cmd_fifo|out_payload[12]~q ),
	.out_payload_13(\clock_crossing_io|cmd_fifo|out_payload[13]~q ),
	.out_payload_14(\clock_crossing_io|cmd_fifo|out_payload[14]~q ),
	.out_payload_15(\clock_crossing_io|cmd_fifo|out_payload[15]~q ),
	.out_payload_16(\clock_crossing_io|cmd_fifo|out_payload[16]~q ),
	.out_payload_17(\clock_crossing_io|cmd_fifo|out_payload[17]~q ),
	.out_payload_18(\clock_crossing_io|cmd_fifo|out_payload[18]~q ),
	.out_payload_19(\clock_crossing_io|cmd_fifo|out_payload[19]~q ),
	.out_payload_20(\clock_crossing_io|cmd_fifo|out_payload[20]~q ),
	.out_payload_0(\clock_crossing_io|rsp_fifo|out_payload[0]~q ),
	.out_payload_1(\clock_crossing_io|rsp_fifo|out_payload[1]~q ),
	.out_payload_2(\clock_crossing_io|rsp_fifo|out_payload[2]~q ),
	.out_payload_3(\clock_crossing_io|rsp_fifo|out_payload[3]~q ),
	.out_payload_4(\clock_crossing_io|rsp_fifo|out_payload[4]~q ),
	.out_payload_51(\clock_crossing_io|rsp_fifo|out_payload[5]~q ),
	.out_payload_61(\clock_crossing_io|rsp_fifo|out_payload[6]~q ),
	.out_payload_71(\clock_crossing_io|rsp_fifo|out_payload[7]~q ),
	.out_payload_81(\clock_crossing_io|rsp_fifo|out_payload[8]~q ),
	.out_payload_91(\clock_crossing_io|rsp_fifo|out_payload[9]~q ),
	.out_payload_101(\clock_crossing_io|rsp_fifo|out_payload[10]~q ),
	.out_payload_111(\clock_crossing_io|rsp_fifo|out_payload[11]~q ),
	.out_payload_121(\clock_crossing_io|rsp_fifo|out_payload[12]~q ),
	.out_payload_131(\clock_crossing_io|rsp_fifo|out_payload[13]~q ),
	.out_payload_141(\clock_crossing_io|rsp_fifo|out_payload[14]~q ),
	.out_payload_151(\clock_crossing_io|rsp_fifo|out_payload[15]~q ),
	.av_readdata_pre_0(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[15]~q ),
	.m0_read1(\mm_interconnect_0|clock_crossing_io_s0_agent|m0_read~2_combout ),
	.m0_write1(\mm_interconnect_0|clock_crossing_io_s0_agent|m0_write~3_combout ),
	.clk_clk(\clk_clk~input_o ));

usb_system_altera_reset_controller_1 rst_controller_001(
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

usb_system_altera_reset_controller rst_controller(
	.wire_pll7_clk_1(\clocks|sd1|wire_pll7_clk[1] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.resetrequest(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_oci_debug|resetrequest~q ),
	.merged_reset(\rst_controller|merged_reset~0_combout ),
	.reset_reset_n(\reset_reset_n~input_o ));

usb_system_altera_irq_clock_crosser irq_synchronizer(
	.r_sync_rst(\rst_controller_002|r_sync_rst~q ),
	.dreg_1(\irq_synchronizer|sync|sync[0].u|dreg[1]~q ),
	.oINT(\cy7c67200_if_0|oINT~q ),
	.clk_clk(\clk_clk~input_o ));

usb_system_usb_system_mm_interconnect_1 mm_interconnect_1(
	.wire_pll7_clk_1(\clocks|sd1|wire_pll7_clk[1] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_valid(\clock_crossing_io|cmd_fifo|out_valid~q ),
	.m0_read(\clock_crossing_io|m0_read~0_combout ),
	.CY7C67200_IF_0_hpi_read(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_read~0_combout ),
	.out_payload_37(\clock_crossing_io|cmd_fifo|out_payload[37]~q ),
	.CY7C67200_IF_0_hpi_write(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_write~0_combout ),
	.waitrequest_reset_override(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|waitrequest_reset_override~q ),
	.av_waitrequest_generated(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_waitrequest_generated~1_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_readdata_pre[15]~q ),
	.oDATA_0(\cy7c67200_if_0|oDATA[0]~q ),
	.oDATA_1(\cy7c67200_if_0|oDATA[1]~q ),
	.oDATA_2(\cy7c67200_if_0|oDATA[2]~q ),
	.oDATA_3(\cy7c67200_if_0|oDATA[3]~q ),
	.oDATA_4(\cy7c67200_if_0|oDATA[4]~q ),
	.oDATA_5(\cy7c67200_if_0|oDATA[5]~q ),
	.oDATA_6(\cy7c67200_if_0|oDATA[6]~q ),
	.oDATA_7(\cy7c67200_if_0|oDATA[7]~q ),
	.oDATA_8(\cy7c67200_if_0|oDATA[8]~q ),
	.oDATA_9(\cy7c67200_if_0|oDATA[9]~q ),
	.oDATA_10(\cy7c67200_if_0|oDATA[10]~q ),
	.oDATA_11(\cy7c67200_if_0|oDATA[11]~q ),
	.oDATA_12(\cy7c67200_if_0|oDATA[12]~q ),
	.oDATA_13(\cy7c67200_if_0|oDATA[13]~q ),
	.oDATA_14(\cy7c67200_if_0|oDATA[14]~q ),
	.oDATA_15(\cy7c67200_if_0|oDATA[15]~q ),
	.av_begintransfer(\mm_interconnect_1|cy7c67200_if_0_hpi_translator|av_begintransfer~2_combout ));

usb_system_altera_reset_controller_3 rst_controller_003(
	.wire_pll7_clk_0(\clocks|sd1|wire_pll7_clk[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_003|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.merged_reset(\rst_controller|merged_reset~0_combout ));

usb_system_altera_reset_controller_2 rst_controller_002(
	.r_sync_rst1(\rst_controller_002|r_sync_rst~q ),
	.merged_reset(\rst_controller|merged_reset~0_combout ),
	.r_early_rst1(\rst_controller_002|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller_002|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .lut_mask = 16'h8BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .sum_lutc_input = "datac";

assign \sdram_wire_dq[0]~input_o  = sdram_wire_dq[0];

assign \sdram_wire_dq[1]~input_o  = sdram_wire_dq[1];

assign \sdram_wire_dq[2]~input_o  = sdram_wire_dq[2];

assign \sdram_wire_dq[3]~input_o  = sdram_wire_dq[3];

assign \sdram_wire_dq[4]~input_o  = sdram_wire_dq[4];

assign \sdram_wire_dq[5]~input_o  = sdram_wire_dq[5];

assign \sdram_wire_dq[6]~input_o  = sdram_wire_dq[6];

assign \sdram_wire_dq[7]~input_o  = sdram_wire_dq[7];

assign \sdram_wire_dq[8]~input_o  = sdram_wire_dq[8];

assign \sdram_wire_dq[9]~input_o  = sdram_wire_dq[9];

assign \sdram_wire_dq[10]~input_o  = sdram_wire_dq[10];

assign \sdram_wire_dq[11]~input_o  = sdram_wire_dq[11];

assign \sdram_wire_dq[12]~input_o  = sdram_wire_dq[12];

assign \sdram_wire_dq[13]~input_o  = sdram_wire_dq[13];

assign \sdram_wire_dq[14]~input_o  = sdram_wire_dq[14];

assign \sdram_wire_dq[15]~input_o  = sdram_wire_dq[15];

assign \sdram_wire_dq[16]~input_o  = sdram_wire_dq[16];

assign \sdram_wire_dq[17]~input_o  = sdram_wire_dq[17];

assign \sdram_wire_dq[18]~input_o  = sdram_wire_dq[18];

assign \sdram_wire_dq[19]~input_o  = sdram_wire_dq[19];

assign \sdram_wire_dq[20]~input_o  = sdram_wire_dq[20];

assign \sdram_wire_dq[21]~input_o  = sdram_wire_dq[21];

assign \sdram_wire_dq[22]~input_o  = sdram_wire_dq[22];

assign \sdram_wire_dq[23]~input_o  = sdram_wire_dq[23];

assign \sdram_wire_dq[24]~input_o  = sdram_wire_dq[24];

assign \sdram_wire_dq[25]~input_o  = sdram_wire_dq[25];

assign \sdram_wire_dq[26]~input_o  = sdram_wire_dq[26];

assign \sdram_wire_dq[27]~input_o  = sdram_wire_dq[27];

assign \sdram_wire_dq[28]~input_o  = sdram_wire_dq[28];

assign \sdram_wire_dq[29]~input_o  = sdram_wire_dq[29];

assign \sdram_wire_dq[30]~input_o  = sdram_wire_dq[30];

assign \sdram_wire_dq[31]~input_o  = sdram_wire_dq[31];

assign \usb_DATA[0]~input_o  = usb_DATA[0];

assign \usb_DATA[1]~input_o  = usb_DATA[1];

assign \usb_DATA[2]~input_o  = usb_DATA[2];

assign \usb_DATA[3]~input_o  = usb_DATA[3];

assign \usb_DATA[4]~input_o  = usb_DATA[4];

assign \usb_DATA[5]~input_o  = usb_DATA[5];

assign \usb_DATA[6]~input_o  = usb_DATA[6];

assign \usb_DATA[7]~input_o  = usb_DATA[7];

assign \usb_DATA[8]~input_o  = usb_DATA[8];

assign \usb_DATA[9]~input_o  = usb_DATA[9];

assign \usb_DATA[10]~input_o  = usb_DATA[10];

assign \usb_DATA[11]~input_o  = usb_DATA[11];

assign \usb_DATA[12]~input_o  = usb_DATA[12];

assign \usb_DATA[13]~input_o  = usb_DATA[13];

assign \usb_DATA[14]~input_o  = usb_DATA[14];

assign \usb_DATA[15]~input_o  = usb_DATA[15];

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \all_switches_wire_export[0]~input_o  = all_switches_wire_export[0];

assign \all_switches_wire_export[1]~input_o  = all_switches_wire_export[1];

assign \all_switches_wire_export[2]~input_o  = all_switches_wire_export[2];

assign \all_switches_wire_export[3]~input_o  = all_switches_wire_export[3];

assign \all_switches_wire_export[4]~input_o  = all_switches_wire_export[4];

assign \all_switches_wire_export[5]~input_o  = all_switches_wire_export[5];

assign \all_switches_wire_export[6]~input_o  = all_switches_wire_export[6];

assign \all_switches_wire_export[7]~input_o  = all_switches_wire_export[7];

assign \all_switches_wire_export[8]~input_o  = all_switches_wire_export[8];

assign \all_switches_wire_export[9]~input_o  = all_switches_wire_export[9];

assign \all_switches_wire_export[10]~input_o  = all_switches_wire_export[10];

assign \all_switches_wire_export[11]~input_o  = all_switches_wire_export[11];

assign \all_switches_wire_export[12]~input_o  = all_switches_wire_export[12];

assign \all_switches_wire_export[13]~input_o  = all_switches_wire_export[13];

assign \all_switches_wire_export[14]~input_o  = all_switches_wire_export[14];

assign \all_switches_wire_export[15]~input_o  = all_switches_wire_export[15];

assign \all_switches_wire_export[16]~input_o  = all_switches_wire_export[16];

assign \all_switches_wire_export[17]~input_o  = all_switches_wire_export[17];

assign \usb_INT~input_o  = usb_INT;

assign keycode_export[0] = \keycode|data_out[0]~q ;

assign keycode_export[1] = \keycode|data_out[1]~q ;

assign keycode_export[2] = \keycode|data_out[2]~q ;

assign keycode_export[3] = \keycode|data_out[3]~q ;

assign keycode_export[4] = \keycode|data_out[4]~q ;

assign keycode_export[5] = \keycode|data_out[5]~q ;

assign keycode_export[6] = \keycode|data_out[6]~q ;

assign keycode_export[7] = \keycode|data_out[7]~q ;

assign led_wire_export[0] = \led|data_out[0]~q ;

assign led_wire_export[1] = \led|data_out[1]~q ;

assign led_wire_export[2] = \led|data_out[2]~q ;

assign led_wire_export[3] = \led|data_out[3]~q ;

assign led_wire_export[4] = \led|data_out[4]~q ;

assign led_wire_export[5] = \led|data_out[5]~q ;

assign led_wire_export[6] = \led|data_out[6]~q ;

assign led_wire_export[7] = \led|data_out[7]~q ;

assign red_leds_wire_export[0] = \red_leds|data_out[0]~q ;

assign red_leds_wire_export[1] = \red_leds|data_out[1]~q ;

assign red_leds_wire_export[2] = \red_leds|data_out[2]~q ;

assign red_leds_wire_export[3] = \red_leds|data_out[3]~q ;

assign red_leds_wire_export[4] = \red_leds|data_out[4]~q ;

assign red_leds_wire_export[5] = \red_leds|data_out[5]~q ;

assign red_leds_wire_export[6] = \red_leds|data_out[6]~q ;

assign red_leds_wire_export[7] = \red_leds|data_out[7]~q ;

assign red_leds_wire_export[8] = \red_leds|data_out[8]~q ;

assign red_leds_wire_export[9] = \red_leds|data_out[9]~q ;

assign red_leds_wire_export[10] = \red_leds|data_out[10]~q ;

assign red_leds_wire_export[11] = \red_leds|data_out[11]~q ;

assign red_leds_wire_export[12] = \red_leds|data_out[12]~q ;

assign red_leds_wire_export[13] = \red_leds|data_out[13]~q ;

assign red_leds_wire_export[14] = \red_leds|data_out[14]~q ;

assign red_leds_wire_export[15] = \red_leds|data_out[15]~q ;

assign red_leds_wire_export[16] = \red_leds|data_out[16]~q ;

assign red_leds_wire_export[17] = \red_leds|data_out[17]~q ;

assign sdram_out_clk_clk = \clocks|sd1|wire_pll7_clk[0] ;

assign sdram_wire_addr[0] = \sdram|m_addr[0]~q ;

assign sdram_wire_addr[1] = \sdram|m_addr[1]~q ;

assign sdram_wire_addr[2] = \sdram|m_addr[2]~q ;

assign sdram_wire_addr[3] = \sdram|m_addr[3]~q ;

assign sdram_wire_addr[4] = \sdram|m_addr[4]~q ;

assign sdram_wire_addr[5] = \sdram|m_addr[5]~q ;

assign sdram_wire_addr[6] = \sdram|m_addr[6]~q ;

assign sdram_wire_addr[7] = \sdram|m_addr[7]~q ;

assign sdram_wire_addr[8] = \sdram|m_addr[8]~q ;

assign sdram_wire_addr[9] = \sdram|m_addr[9]~q ;

assign sdram_wire_addr[10] = \sdram|m_addr[10]~q ;

assign sdram_wire_addr[11] = \sdram|m_addr[11]~q ;

assign sdram_wire_addr[12] = \sdram|m_addr[12]~q ;

assign sdram_wire_ba[0] = \sdram|m_bank[0]~q ;

assign sdram_wire_ba[1] = \sdram|m_bank[1]~q ;

assign sdram_wire_cas_n = ~ \sdram|m_cmd[1]~q ;

assign sdram_wire_cke = vcc;

assign sdram_wire_cs_n = ~ \sdram|m_cmd[3]~q ;

assign sdram_wire_dqm[0] = \sdram|m_dqm[0]~q ;

assign sdram_wire_dqm[1] = \sdram|m_dqm[1]~q ;

assign sdram_wire_dqm[2] = \sdram|m_dqm[2]~q ;

assign sdram_wire_dqm[3] = \sdram|m_dqm[3]~q ;

assign sdram_wire_ras_n = ~ \sdram|m_cmd[2]~q ;

assign sdram_wire_we_n = ~ \sdram|m_cmd[0]~q ;

assign usb_ADDR[0] = \cy7c67200_if_0|HPI_ADDR[0]~q ;

assign usb_ADDR[1] = \cy7c67200_if_0|HPI_ADDR[1]~q ;

assign usb_RD_N = ~ \cy7c67200_if_0|HPI_RD_N~q ;

assign usb_WR_N = ~ \cy7c67200_if_0|HPI_WR_N~q ;

assign usb_CS_N = ~ \cy7c67200_if_0|HPI_CS_N~q ;

assign usb_RST_N = \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;

assign usb_out_clk_clk = \clocks|sd1|wire_pll7_clk[1] ;

cycloneive_io_obuf \sdram_wire_dq[0]~output (
	.i(\sdram|m_data[0]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[0]),
	.obar());
defparam \sdram_wire_dq[0]~output .bus_hold = "false";
defparam \sdram_wire_dq[0]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[1]~output (
	.i(\sdram|m_data[1]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[1]),
	.obar());
defparam \sdram_wire_dq[1]~output .bus_hold = "false";
defparam \sdram_wire_dq[1]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[2]~output (
	.i(\sdram|m_data[2]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[2]),
	.obar());
defparam \sdram_wire_dq[2]~output .bus_hold = "false";
defparam \sdram_wire_dq[2]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[3]~output (
	.i(\sdram|m_data[3]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[3]),
	.obar());
defparam \sdram_wire_dq[3]~output .bus_hold = "false";
defparam \sdram_wire_dq[3]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[4]~output (
	.i(\sdram|m_data[4]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[4]),
	.obar());
defparam \sdram_wire_dq[4]~output .bus_hold = "false";
defparam \sdram_wire_dq[4]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[5]~output (
	.i(\sdram|m_data[5]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[5]),
	.obar());
defparam \sdram_wire_dq[5]~output .bus_hold = "false";
defparam \sdram_wire_dq[5]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[6]~output (
	.i(\sdram|m_data[6]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[6]),
	.obar());
defparam \sdram_wire_dq[6]~output .bus_hold = "false";
defparam \sdram_wire_dq[6]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[7]~output (
	.i(\sdram|m_data[7]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[7]),
	.obar());
defparam \sdram_wire_dq[7]~output .bus_hold = "false";
defparam \sdram_wire_dq[7]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[8]~output (
	.i(\sdram|m_data[8]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[8]),
	.obar());
defparam \sdram_wire_dq[8]~output .bus_hold = "false";
defparam \sdram_wire_dq[8]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[9]~output (
	.i(\sdram|m_data[9]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[9]),
	.obar());
defparam \sdram_wire_dq[9]~output .bus_hold = "false";
defparam \sdram_wire_dq[9]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[10]~output (
	.i(\sdram|m_data[10]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[10]),
	.obar());
defparam \sdram_wire_dq[10]~output .bus_hold = "false";
defparam \sdram_wire_dq[10]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[11]~output (
	.i(\sdram|m_data[11]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[11]),
	.obar());
defparam \sdram_wire_dq[11]~output .bus_hold = "false";
defparam \sdram_wire_dq[11]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[12]~output (
	.i(\sdram|m_data[12]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[12]),
	.obar());
defparam \sdram_wire_dq[12]~output .bus_hold = "false";
defparam \sdram_wire_dq[12]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[13]~output (
	.i(\sdram|m_data[13]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[13]),
	.obar());
defparam \sdram_wire_dq[13]~output .bus_hold = "false";
defparam \sdram_wire_dq[13]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[14]~output (
	.i(\sdram|m_data[14]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[14]),
	.obar());
defparam \sdram_wire_dq[14]~output .bus_hold = "false";
defparam \sdram_wire_dq[14]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[15]~output (
	.i(\sdram|m_data[15]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[15]),
	.obar());
defparam \sdram_wire_dq[15]~output .bus_hold = "false";
defparam \sdram_wire_dq[15]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[16]~output (
	.i(\sdram|m_data[16]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[16]),
	.obar());
defparam \sdram_wire_dq[16]~output .bus_hold = "false";
defparam \sdram_wire_dq[16]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[17]~output (
	.i(\sdram|m_data[17]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[17]),
	.obar());
defparam \sdram_wire_dq[17]~output .bus_hold = "false";
defparam \sdram_wire_dq[17]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[18]~output (
	.i(\sdram|m_data[18]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[18]),
	.obar());
defparam \sdram_wire_dq[18]~output .bus_hold = "false";
defparam \sdram_wire_dq[18]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[19]~output (
	.i(\sdram|m_data[19]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[19]),
	.obar());
defparam \sdram_wire_dq[19]~output .bus_hold = "false";
defparam \sdram_wire_dq[19]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[20]~output (
	.i(\sdram|m_data[20]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[20]),
	.obar());
defparam \sdram_wire_dq[20]~output .bus_hold = "false";
defparam \sdram_wire_dq[20]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[21]~output (
	.i(\sdram|m_data[21]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[21]),
	.obar());
defparam \sdram_wire_dq[21]~output .bus_hold = "false";
defparam \sdram_wire_dq[21]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[22]~output (
	.i(\sdram|m_data[22]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[22]),
	.obar());
defparam \sdram_wire_dq[22]~output .bus_hold = "false";
defparam \sdram_wire_dq[22]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[23]~output (
	.i(\sdram|m_data[23]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[23]),
	.obar());
defparam \sdram_wire_dq[23]~output .bus_hold = "false";
defparam \sdram_wire_dq[23]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[24]~output (
	.i(\sdram|m_data[24]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[24]),
	.obar());
defparam \sdram_wire_dq[24]~output .bus_hold = "false";
defparam \sdram_wire_dq[24]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[25]~output (
	.i(\sdram|m_data[25]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[25]),
	.obar());
defparam \sdram_wire_dq[25]~output .bus_hold = "false";
defparam \sdram_wire_dq[25]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[26]~output (
	.i(\sdram|m_data[26]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[26]),
	.obar());
defparam \sdram_wire_dq[26]~output .bus_hold = "false";
defparam \sdram_wire_dq[26]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[27]~output (
	.i(\sdram|m_data[27]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[27]),
	.obar());
defparam \sdram_wire_dq[27]~output .bus_hold = "false";
defparam \sdram_wire_dq[27]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[28]~output (
	.i(\sdram|m_data[28]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[28]),
	.obar());
defparam \sdram_wire_dq[28]~output .bus_hold = "false";
defparam \sdram_wire_dq[28]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[29]~output (
	.i(\sdram|m_data[29]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[29]),
	.obar());
defparam \sdram_wire_dq[29]~output .bus_hold = "false";
defparam \sdram_wire_dq[29]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[30]~output (
	.i(\sdram|m_data[30]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[30]),
	.obar());
defparam \sdram_wire_dq[30]~output .bus_hold = "false";
defparam \sdram_wire_dq[30]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[31]~output (
	.i(\sdram|m_data[31]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[31]),
	.obar());
defparam \sdram_wire_dq[31]~output .bus_hold = "false";
defparam \sdram_wire_dq[31]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[0]~output (
	.i(\cy7c67200_if_0|TMP_DATA[0]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[0]),
	.obar());
defparam \usb_DATA[0]~output .bus_hold = "false";
defparam \usb_DATA[0]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[1]~output (
	.i(\cy7c67200_if_0|TMP_DATA[1]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[1]),
	.obar());
defparam \usb_DATA[1]~output .bus_hold = "false";
defparam \usb_DATA[1]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[2]~output (
	.i(\cy7c67200_if_0|TMP_DATA[2]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[2]),
	.obar());
defparam \usb_DATA[2]~output .bus_hold = "false";
defparam \usb_DATA[2]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[3]~output (
	.i(\cy7c67200_if_0|TMP_DATA[3]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[3]),
	.obar());
defparam \usb_DATA[3]~output .bus_hold = "false";
defparam \usb_DATA[3]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[4]~output (
	.i(\cy7c67200_if_0|TMP_DATA[4]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[4]),
	.obar());
defparam \usb_DATA[4]~output .bus_hold = "false";
defparam \usb_DATA[4]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[5]~output (
	.i(\cy7c67200_if_0|TMP_DATA[5]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[5]),
	.obar());
defparam \usb_DATA[5]~output .bus_hold = "false";
defparam \usb_DATA[5]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[6]~output (
	.i(\cy7c67200_if_0|TMP_DATA[6]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[6]),
	.obar());
defparam \usb_DATA[6]~output .bus_hold = "false";
defparam \usb_DATA[6]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[7]~output (
	.i(\cy7c67200_if_0|TMP_DATA[7]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[7]),
	.obar());
defparam \usb_DATA[7]~output .bus_hold = "false";
defparam \usb_DATA[7]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[8]~output (
	.i(\cy7c67200_if_0|TMP_DATA[8]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[8]),
	.obar());
defparam \usb_DATA[8]~output .bus_hold = "false";
defparam \usb_DATA[8]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[9]~output (
	.i(\cy7c67200_if_0|TMP_DATA[9]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[9]),
	.obar());
defparam \usb_DATA[9]~output .bus_hold = "false";
defparam \usb_DATA[9]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[10]~output (
	.i(\cy7c67200_if_0|TMP_DATA[10]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[10]),
	.obar());
defparam \usb_DATA[10]~output .bus_hold = "false";
defparam \usb_DATA[10]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[11]~output (
	.i(\cy7c67200_if_0|TMP_DATA[11]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[11]),
	.obar());
defparam \usb_DATA[11]~output .bus_hold = "false";
defparam \usb_DATA[11]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[12]~output (
	.i(\cy7c67200_if_0|TMP_DATA[12]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[12]),
	.obar());
defparam \usb_DATA[12]~output .bus_hold = "false";
defparam \usb_DATA[12]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[13]~output (
	.i(\cy7c67200_if_0|TMP_DATA[13]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[13]),
	.obar());
defparam \usb_DATA[13]~output .bus_hold = "false";
defparam \usb_DATA[13]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[14]~output (
	.i(\cy7c67200_if_0|TMP_DATA[14]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[14]),
	.obar());
defparam \usb_DATA[14]~output .bus_hold = "false";
defparam \usb_DATA[14]~output .open_drain_output = "false";

cycloneive_io_obuf \usb_DATA[15]~output (
	.i(\cy7c67200_if_0|TMP_DATA[15]~q ),
	.oe(\cy7c67200_if_0|HPI_WR_N~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(usb_DATA[15]),
	.obar());
defparam \usb_DATA[15]~output .bus_hold = "false";
defparam \usb_DATA[15]~output .open_drain_output = "false";

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~10 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~10 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 .lut_mask = 16'hCF5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0 (
	.dataa(\~GND~combout ),
	.datab(\rst_controller_002|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 16'hBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .lut_mask = 16'h9696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2_combout ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .lut_mask = 16'hBEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14 .lut_mask = 16'hDDF5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0_combout ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8 .lut_mask = 16'hFFDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'h7777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .lut_mask = 16'hBFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .lut_mask = 16'hFF6F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .lut_mask = 16'hFFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 (
	.dataa(\cpu|cpu|the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\jtag_uart|usb_system_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_mm_clock_crossing_bridge (
	wire_pll7_clk_1,
	W_alu_result_2,
	W_alu_result_3,
	m0_reset,
	d_writedata_0,
	r_sync_rst,
	d_write,
	write_accepted,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	out_payload_42,
	out_payload_43,
	out_valid,
	m0_read,
	out_payload_37,
	sink_in_reset,
	d_read,
	read_accepted,
	out_valid1,
	full,
	s0_cmd_valid1,
	waitrequest_reset_override,
	av_waitrequest_generated,
	m0_write,
	read_latency_shift_reg_0,
	out_payload_5,
	out_payload_6,
	out_payload_7,
	out_payload_8,
	out_payload_9,
	out_payload_10,
	out_payload_11,
	out_payload_12,
	out_payload_13,
	out_payload_14,
	out_payload_15,
	out_payload_16,
	out_payload_17,
	out_payload_18,
	out_payload_19,
	out_payload_20,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_51,
	out_payload_61,
	out_payload_71,
	out_payload_81,
	out_payload_91,
	out_payload_101,
	out_payload_111,
	out_payload_121,
	out_payload_131,
	out_payload_141,
	out_payload_151,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	m0_read1,
	m0_write1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	m0_reset;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_write;
input 	write_accepted;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
output 	out_payload_42;
output 	out_payload_43;
output 	out_valid;
output 	m0_read;
output 	out_payload_37;
output 	sink_in_reset;
input 	d_read;
input 	read_accepted;
output 	out_valid1;
output 	full;
output 	s0_cmd_valid1;
input 	waitrequest_reset_override;
input 	av_waitrequest_generated;
input 	m0_write;
input 	read_latency_shift_reg_0;
output 	out_payload_5;
output 	out_payload_6;
output 	out_payload_7;
output 	out_payload_8;
output 	out_payload_9;
output 	out_payload_10;
output 	out_payload_11;
output 	out_payload_12;
output 	out_payload_13;
output 	out_payload_14;
output 	out_payload_15;
output 	out_payload_16;
output 	out_payload_17;
output 	out_payload_18;
output 	out_payload_19;
output 	out_payload_20;
output 	out_payload_0;
output 	out_payload_1;
output 	out_payload_2;
output 	out_payload_3;
output 	out_payload_4;
output 	out_payload_51;
output 	out_payload_61;
output 	out_payload_71;
output 	out_payload_81;
output 	out_payload_91;
output 	out_payload_101;
output 	out_payload_111;
output 	out_payload_121;
output 	out_payload_131;
output 	out_payload_141;
output 	out_payload_151;
input 	av_readdata_pre_0;
input 	av_readdata_pre_1;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_7;
input 	av_readdata_pre_8;
input 	av_readdata_pre_9;
input 	av_readdata_pre_10;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	m0_read1;
input 	m0_write1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rsp_fifo|in_space_avail[8]~q ;
wire \rsp_fifo|in_space_avail[7]~q ;
wire \rsp_fifo|in_space_avail[6]~q ;
wire \rsp_fifo|in_space_avail[5]~q ;
wire \rsp_fifo|in_space_avail[4]~q ;
wire \rsp_fifo|in_space_avail[3]~q ;
wire \rsp_fifo|in_space_avail[2]~q ;
wire \rsp_fifo|in_space_avail[1]~q ;
wire \rsp_fifo|in_space_avail[0]~q ;
wire \cmd_fifo|out_payload[38]~q ;
wire \old_read~0_combout ;
wire \old_read~q ;
wire \pending_read_count[0]~9_combout ;
wire \pending_read_count[1]~27_combout ;
wire \pending_read_count[0]~q ;
wire \pending_read_count[0]~10 ;
wire \pending_read_count[1]~11_combout ;
wire \pending_read_count[1]~q ;
wire \pending_read_count[1]~12 ;
wire \pending_read_count[2]~13_combout ;
wire \pending_read_count[2]~q ;
wire \pending_read_count[2]~14 ;
wire \pending_read_count[3]~15_combout ;
wire \pending_read_count[3]~q ;
wire \pending_read_count[3]~16 ;
wire \pending_read_count[4]~17_combout ;
wire \pending_read_count[4]~q ;
wire \pending_read_count[4]~18 ;
wire \pending_read_count[5]~19_combout ;
wire \pending_read_count[5]~q ;
wire \pending_read_count[5]~20 ;
wire \pending_read_count[6]~21_combout ;
wire \pending_read_count[6]~q ;
wire \pending_read_count[6]~22 ;
wire \pending_read_count[7]~23_combout ;
wire \pending_read_count[7]~q ;
wire \pending_read_count[7]~24 ;
wire \pending_read_count[8]~25_combout ;
wire \pending_read_count[8]~q ;
wire \Add2~1 ;
wire \Add2~3 ;
wire \Add2~5 ;
wire \Add2~7 ;
wire \Add2~9 ;
wire \Add2~11 ;
wire \Add2~12_combout ;
wire \Add2~10_combout ;
wire \Add2~8_combout ;
wire \Add2~6_combout ;
wire \Add2~4_combout ;
wire \Add2~2_combout ;
wire \Add2~0_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~16_combout ;
wire \Add2~13 ;
wire \Add2~14_combout ;
wire \LessThan0~18_combout ;
wire \stop_cmd_r~q ;


usb_system_altera_avalon_dc_fifo_1 rsp_fifo(
	.wire_pll7_clk_1(wire_pll7_clk_1),
	.in_space_avail_8(\rsp_fifo|in_space_avail[8]~q ),
	.in_space_avail_7(\rsp_fifo|in_space_avail[7]~q ),
	.in_space_avail_6(\rsp_fifo|in_space_avail[6]~q ),
	.in_space_avail_5(\rsp_fifo|in_space_avail[5]~q ),
	.in_space_avail_4(\rsp_fifo|in_space_avail[4]~q ),
	.in_space_avail_3(\rsp_fifo|in_space_avail[3]~q ),
	.in_space_avail_2(\rsp_fifo|in_space_avail[2]~q ),
	.in_space_avail_1(\rsp_fifo|in_space_avail[1]~q ),
	.in_space_avail_0(\rsp_fifo|in_space_avail[0]~q ),
	.altera_reset_synchronizer_int_chain_out(m0_reset),
	.r_sync_rst(r_sync_rst),
	.out_valid1(out_valid1),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.out_payload_0(out_payload_0),
	.out_payload_1(out_payload_1),
	.out_payload_2(out_payload_2),
	.out_payload_3(out_payload_3),
	.out_payload_4(out_payload_4),
	.out_payload_5(out_payload_51),
	.out_payload_6(out_payload_61),
	.out_payload_7(out_payload_71),
	.out_payload_8(out_payload_81),
	.out_payload_9(out_payload_91),
	.out_payload_10(out_payload_101),
	.out_payload_11(out_payload_111),
	.out_payload_12(out_payload_121),
	.out_payload_13(out_payload_131),
	.out_payload_14(out_payload_141),
	.out_payload_15(out_payload_151),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.clk_clk(clk_clk));

usb_system_altera_avalon_dc_fifo cmd_fifo(
	.wire_pll7_clk_1(wire_pll7_clk_1),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.altera_reset_synchronizer_int_chain_out(m0_reset),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.out_payload_42(out_payload_42),
	.out_payload_43(out_payload_43),
	.out_valid1(out_valid),
	.out_payload_38(\cmd_fifo|out_payload[38]~q ),
	.old_read(\old_read~q ),
	.stop_cmd_r(\stop_cmd_r~q ),
	.out_payload_37(out_payload_37),
	.sink_in_reset1(sink_in_reset),
	.full1(full),
	.s0_cmd_valid(s0_cmd_valid1),
	.waitrequest_reset_override(waitrequest_reset_override),
	.av_waitrequest_generated(av_waitrequest_generated),
	.m0_write(m0_write),
	.out_payload_5(out_payload_5),
	.out_payload_6(out_payload_6),
	.out_payload_7(out_payload_7),
	.out_payload_8(out_payload_8),
	.out_payload_9(out_payload_9),
	.out_payload_10(out_payload_10),
	.out_payload_11(out_payload_11),
	.out_payload_12(out_payload_12),
	.out_payload_13(out_payload_13),
	.out_payload_14(out_payload_14),
	.out_payload_15(out_payload_15),
	.out_payload_16(out_payload_16),
	.out_payload_17(out_payload_17),
	.out_payload_18(out_payload_18),
	.out_payload_19(out_payload_19),
	.out_payload_20(out_payload_20),
	.m0_read(m0_read1),
	.m0_write1(m0_write1),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \m0_read~0 (
	.dataa(out_valid),
	.datab(\cmd_fifo|out_payload[38]~q ),
	.datac(\old_read~q ),
	.datad(\stop_cmd_r~q ),
	.cin(gnd),
	.combout(m0_read),
	.cout());
defparam \m0_read~0 .lut_mask = 16'hFEFF;
defparam \m0_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb s0_cmd_valid(
	.dataa(d_write),
	.datab(d_read),
	.datac(write_accepted),
	.datad(read_accepted),
	.cin(gnd),
	.combout(s0_cmd_valid1),
	.cout());
defparam s0_cmd_valid.lut_mask = 16'hEFFF;
defparam s0_cmd_valid.sum_lutc_input = "datac";

cycloneive_lcell_comb \old_read~0 (
	.dataa(m0_read),
	.datab(av_waitrequest_generated),
	.datac(gnd),
	.datad(waitrequest_reset_override),
	.cin(gnd),
	.combout(\old_read~0_combout ),
	.cout());
defparam \old_read~0 .lut_mask = 16'hEEFF;
defparam \old_read~0 .sum_lutc_input = "datac";

dffeas old_read(
	.clk(wire_pll7_clk_1),
	.d(\old_read~0_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\old_read~q ),
	.prn(vcc));
defparam old_read.is_wysiwyg = "true";
defparam old_read.power_up = "low";

cycloneive_lcell_comb \pending_read_count[0]~9 (
	.dataa(\pending_read_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\pending_read_count[0]~9_combout ),
	.cout(\pending_read_count[0]~10 ));
defparam \pending_read_count[0]~9 .lut_mask = 16'h55AA;
defparam \pending_read_count[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending_read_count[1]~27 (
	.dataa(m0_read),
	.datab(waitrequest_reset_override),
	.datac(av_waitrequest_generated),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\pending_read_count[1]~27_combout ),
	.cout());
defparam \pending_read_count[1]~27 .lut_mask = 16'h6996;
defparam \pending_read_count[1]~27 .sum_lutc_input = "datac";

dffeas \pending_read_count[0] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[0]~9_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[0]~q ),
	.prn(vcc));
defparam \pending_read_count[0] .is_wysiwyg = "true";
defparam \pending_read_count[0] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[1]~11 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[0]~10 ),
	.combout(\pending_read_count[1]~11_combout ),
	.cout(\pending_read_count[1]~12 ));
defparam \pending_read_count[1]~11 .lut_mask = 16'h967F;
defparam \pending_read_count[1]~11 .sum_lutc_input = "cin";

dffeas \pending_read_count[1] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[1]~11_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[1]~q ),
	.prn(vcc));
defparam \pending_read_count[1] .is_wysiwyg = "true";
defparam \pending_read_count[1] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[2]~13 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[1]~12 ),
	.combout(\pending_read_count[2]~13_combout ),
	.cout(\pending_read_count[2]~14 ));
defparam \pending_read_count[2]~13 .lut_mask = 16'h96EF;
defparam \pending_read_count[2]~13 .sum_lutc_input = "cin";

dffeas \pending_read_count[2] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[2]~13_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[2]~q ),
	.prn(vcc));
defparam \pending_read_count[2] .is_wysiwyg = "true";
defparam \pending_read_count[2] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[3]~15 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[2]~14 ),
	.combout(\pending_read_count[3]~15_combout ),
	.cout(\pending_read_count[3]~16 ));
defparam \pending_read_count[3]~15 .lut_mask = 16'h967F;
defparam \pending_read_count[3]~15 .sum_lutc_input = "cin";

dffeas \pending_read_count[3] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[3]~15_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[3]~q ),
	.prn(vcc));
defparam \pending_read_count[3] .is_wysiwyg = "true";
defparam \pending_read_count[3] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[4]~17 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[3]~16 ),
	.combout(\pending_read_count[4]~17_combout ),
	.cout(\pending_read_count[4]~18 ));
defparam \pending_read_count[4]~17 .lut_mask = 16'h96EF;
defparam \pending_read_count[4]~17 .sum_lutc_input = "cin";

dffeas \pending_read_count[4] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[4]~17_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[4]~q ),
	.prn(vcc));
defparam \pending_read_count[4] .is_wysiwyg = "true";
defparam \pending_read_count[4] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[5]~19 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[4]~18 ),
	.combout(\pending_read_count[5]~19_combout ),
	.cout(\pending_read_count[5]~20 ));
defparam \pending_read_count[5]~19 .lut_mask = 16'h967F;
defparam \pending_read_count[5]~19 .sum_lutc_input = "cin";

dffeas \pending_read_count[5] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[5]~19_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[5]~q ),
	.prn(vcc));
defparam \pending_read_count[5] .is_wysiwyg = "true";
defparam \pending_read_count[5] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[6]~21 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[5]~20 ),
	.combout(\pending_read_count[6]~21_combout ),
	.cout(\pending_read_count[6]~22 ));
defparam \pending_read_count[6]~21 .lut_mask = 16'h96EF;
defparam \pending_read_count[6]~21 .sum_lutc_input = "cin";

dffeas \pending_read_count[6] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[6]~21_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[6]~q ),
	.prn(vcc));
defparam \pending_read_count[6] .is_wysiwyg = "true";
defparam \pending_read_count[6] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[7]~23 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\pending_read_count[6]~22 ),
	.combout(\pending_read_count[7]~23_combout ),
	.cout(\pending_read_count[7]~24 ));
defparam \pending_read_count[7]~23 .lut_mask = 16'h967F;
defparam \pending_read_count[7]~23 .sum_lutc_input = "cin";

dffeas \pending_read_count[7] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[7]~23_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[7]~q ),
	.prn(vcc));
defparam \pending_read_count[7] .is_wysiwyg = "true";
defparam \pending_read_count[7] .power_up = "low";

cycloneive_lcell_comb \pending_read_count[8]~25 (
	.dataa(read_latency_shift_reg_0),
	.datab(\pending_read_count[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\pending_read_count[7]~24 ),
	.combout(\pending_read_count[8]~25_combout ),
	.cout());
defparam \pending_read_count[8]~25 .lut_mask = 16'h9696;
defparam \pending_read_count[8]~25 .sum_lutc_input = "cin";

dffeas \pending_read_count[8] (
	.clk(wire_pll7_clk_1),
	.d(\pending_read_count[8]~25_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_read_count[1]~27_combout ),
	.q(\pending_read_count[8]~q ),
	.prn(vcc));
defparam \pending_read_count[8] .is_wysiwyg = "true";
defparam \pending_read_count[8] .power_up = "low";

cycloneive_lcell_comb \Add2~0 (
	.dataa(\pending_read_count[1]~q ),
	.datab(\pending_read_count[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h66EE;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add2~2 (
	.dataa(\pending_read_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'h5A5F;
defparam \Add2~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~4 (
	.dataa(\pending_read_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h5AAF;
defparam \Add2~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~6 (
	.dataa(\pending_read_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'h5A5F;
defparam \Add2~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~8 (
	.dataa(\pending_read_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
defparam \Add2~8 .lut_mask = 16'h5AAF;
defparam \Add2~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~10 (
	.dataa(\pending_read_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
defparam \Add2~10 .lut_mask = 16'h5A5F;
defparam \Add2~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~12 (
	.dataa(\pending_read_count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
defparam \Add2~12 .lut_mask = 16'h5AAF;
defparam \Add2~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\rsp_fifo|in_space_avail[0]~q ),
	.datab(\pending_read_count[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
defparam \LessThan0~1 .lut_mask = 16'h00DD;
defparam \LessThan0~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~3 (
	.dataa(\rsp_fifo|in_space_avail[1]~q ),
	.datab(\pending_read_count[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
defparam \LessThan0~3 .lut_mask = 16'h00EF;
defparam \LessThan0~3 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~5 (
	.dataa(\rsp_fifo|in_space_avail[2]~q ),
	.datab(\Add2~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
defparam \LessThan0~5 .lut_mask = 16'h00DF;
defparam \LessThan0~5 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~7 (
	.dataa(\rsp_fifo|in_space_avail[3]~q ),
	.datab(\Add2~2_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
defparam \LessThan0~7 .lut_mask = 16'h00BF;
defparam \LessThan0~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~9 (
	.dataa(\rsp_fifo|in_space_avail[4]~q ),
	.datab(\Add2~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
defparam \LessThan0~9 .lut_mask = 16'h00DF;
defparam \LessThan0~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~11 (
	.dataa(\rsp_fifo|in_space_avail[5]~q ),
	.datab(\Add2~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
defparam \LessThan0~11 .lut_mask = 16'h00BF;
defparam \LessThan0~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~13 (
	.dataa(\rsp_fifo|in_space_avail[6]~q ),
	.datab(\Add2~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
defparam \LessThan0~13 .lut_mask = 16'h00DF;
defparam \LessThan0~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~15 (
	.dataa(\rsp_fifo|in_space_avail[7]~q ),
	.datab(\Add2~10_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
defparam \LessThan0~15 .lut_mask = 16'h00BF;
defparam \LessThan0~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~16 (
	.dataa(\rsp_fifo|in_space_avail[8]~q ),
	.datab(\Add2~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan0~15_cout ),
	.combout(\LessThan0~16_combout ),
	.cout());
defparam \LessThan0~16 .lut_mask = 16'hEFEF;
defparam \LessThan0~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout());
defparam \Add2~14 .lut_mask = 16'hF0F0;
defparam \Add2~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan0~18 (
	.dataa(\LessThan0~16_combout ),
	.datab(\Add2~14_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan0~18_combout ),
	.cout());
defparam \LessThan0~18 .lut_mask = 16'hEEEE;
defparam \LessThan0~18 .sum_lutc_input = "datac";

dffeas stop_cmd_r(
	.clk(wire_pll7_clk_1),
	.d(\LessThan0~18_combout ),
	.asdata(vcc),
	.clrn(m0_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stop_cmd_r~q ),
	.prn(vcc));
defparam stop_cmd_r.is_wysiwyg = "true";
defparam stop_cmd_r.power_up = "low";

endmodule

module usb_system_altera_avalon_dc_fifo (
	wire_pll7_clk_1,
	W_alu_result_2,
	W_alu_result_3,
	altera_reset_synchronizer_int_chain_out,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	out_payload_42,
	out_payload_43,
	out_valid1,
	out_payload_38,
	old_read,
	stop_cmd_r,
	out_payload_37,
	sink_in_reset1,
	full1,
	s0_cmd_valid,
	waitrequest_reset_override,
	av_waitrequest_generated,
	m0_write,
	out_payload_5,
	out_payload_6,
	out_payload_7,
	out_payload_8,
	out_payload_9,
	out_payload_10,
	out_payload_11,
	out_payload_12,
	out_payload_13,
	out_payload_14,
	out_payload_15,
	out_payload_16,
	out_payload_17,
	out_payload_18,
	out_payload_19,
	out_payload_20,
	m0_read,
	m0_write1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	altera_reset_synchronizer_int_chain_out;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
output 	out_payload_42;
output 	out_payload_43;
output 	out_valid1;
output 	out_payload_38;
input 	old_read;
input 	stop_cmd_r;
output 	out_payload_37;
output 	sink_in_reset1;
output 	full1;
input 	s0_cmd_valid;
input 	waitrequest_reset_override;
input 	av_waitrequest_generated;
input 	m0_write;
output 	out_payload_5;
output 	out_payload_6;
output 	out_payload_7;
output 	out_payload_8;
output 	out_payload_9;
output 	out_payload_10;
output 	out_payload_11;
output 	out_payload_12;
output 	out_payload_13;
output 	out_payload_14;
output 	out_payload_15;
output 	out_payload_16;
output 	out_payload_17;
output 	out_payload_18;
output 	out_payload_19;
output 	out_payload_20;
input 	m0_read;
input 	m0_write1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_crosser|sync[1].u|dreg[1]~q ;
wire \read_crosser|sync[2].u|dreg[1]~q ;
wire \read_crosser|sync[3].u|dreg[1]~q ;
wire \read_crosser|sync[4].u|dreg[1]~q ;
wire \read_crosser|sync[5].u|dreg[1]~q ;
wire \read_crosser|sync[0].u|dreg[1]~q ;
wire \write_crosser|sync[1].u|dreg[1]~q ;
wire \write_crosser|sync[2].u|dreg[1]~q ;
wire \write_crosser|sync[3].u|dreg[1]~q ;
wire \write_crosser|sync[4].u|dreg[1]~q ;
wire \write_crosser|sync[5].u|dreg[1]~q ;
wire \write_crosser|sync[0].u|dreg[1]~q ;
wire \out_rd_ptr_gray[1]~q ;
wire \out_rd_ptr_gray[2]~q ;
wire \out_rd_ptr_gray[3]~q ;
wire \out_rd_ptr_gray[4]~q ;
wire \out_rd_ptr_gray[5]~q ;
wire \out_rd_ptr_gray[0]~q ;
wire \in_wr_ptr_gray[1]~q ;
wire \in_wr_ptr_gray[2]~q ;
wire \in_wr_ptr_gray[3]~q ;
wire \in_wr_ptr_gray[4]~q ;
wire \in_wr_ptr_gray[5]~q ;
wire \in_wr_ptr_gray[0]~q ;
wire \bin2gray~0_combout ;
wire \bin2gray~1_combout ;
wire \bin2gray~2_combout ;
wire \bin2gray~3_combout ;
wire \bin2gray~4_combout ;
wire \bin2gray~5_combout ;
wire \bin2gray~6_combout ;
wire \bin2gray~7_combout ;
wire \bin2gray~8_combout ;
wire \bin2gray~9_combout ;
wire \next_in_wr_ptr~0_combout ;
wire \Add0~0_combout ;
wire \in_wr_ptr[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \in_wr_ptr[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \in_wr_ptr[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \in_wr_ptr[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \in_wr_ptr[4]~q ;
wire \out_rd_ptr[0]~q ;
wire \internal_out_ready~0_combout ;
wire \internal_out_ready~1_combout ;
wire \out_rd_ptr[1]~q ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \out_rd_ptr[4]~q ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \out_rd_ptr[2]~q ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \out_rd_ptr[3]~q ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \out_rd_ptr[5]~q ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Equal0~6_combout ;
wire \empty~q ;
wire \next_out_rd_ptr~0_combout ;
wire \Add1~0_combout ;
wire \mem_rtl_0|auto_generated|ram_block1a18~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a19~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a17~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a16~portbdataout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \full~0_combout ;
wire \in_wr_ptr[5]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \full~1_combout ;
wire \Equal1~2_combout ;
wire \Equal1~3_combout ;
wire \full~2_combout ;
wire \mem_rtl_0|auto_generated|ram_block1a0~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a1~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a2~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a3~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a4~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a5~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a6~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a7~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a8~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a9~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a10~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a11~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a12~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a13~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a14~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a15~portbdataout ;

wire [143:0] \mem_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ;

assign \mem_rtl_0|auto_generated|ram_block1a18~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a19~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a17~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a16~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a0~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a1~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a2~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a3~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a4~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a5~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a6~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a7~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a8~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a9~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a10~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a11~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a12~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a13~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a14~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a15~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus [0];

usb_system_altera_dcfifo_synchronizer_bundle read_crosser(
	.r_sync_rst(r_sync_rst),
	.dreg_1(\read_crosser|sync[1].u|dreg[1]~q ),
	.dreg_11(\read_crosser|sync[2].u|dreg[1]~q ),
	.dreg_12(\read_crosser|sync[3].u|dreg[1]~q ),
	.dreg_13(\read_crosser|sync[4].u|dreg[1]~q ),
	.dreg_14(\read_crosser|sync[5].u|dreg[1]~q ),
	.dreg_15(\read_crosser|sync[0].u|dreg[1]~q ),
	.out_rd_ptr_gray_1(\out_rd_ptr_gray[1]~q ),
	.out_rd_ptr_gray_2(\out_rd_ptr_gray[2]~q ),
	.out_rd_ptr_gray_3(\out_rd_ptr_gray[3]~q ),
	.out_rd_ptr_gray_4(\out_rd_ptr_gray[4]~q ),
	.out_rd_ptr_gray_5(\out_rd_ptr_gray[5]~q ),
	.out_rd_ptr_gray_0(\out_rd_ptr_gray[0]~q ),
	.clk_clk(clk_clk));

usb_system_altera_dcfifo_synchronizer_bundle_1 write_crosser(
	.wire_pll7_clk_1(wire_pll7_clk_1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.dreg_1(\write_crosser|sync[1].u|dreg[1]~q ),
	.dreg_11(\write_crosser|sync[2].u|dreg[1]~q ),
	.dreg_12(\write_crosser|sync[3].u|dreg[1]~q ),
	.dreg_13(\write_crosser|sync[4].u|dreg[1]~q ),
	.dreg_14(\write_crosser|sync[5].u|dreg[1]~q ),
	.dreg_15(\write_crosser|sync[0].u|dreg[1]~q ),
	.in_wr_ptr_gray_1(\in_wr_ptr_gray[1]~q ),
	.in_wr_ptr_gray_2(\in_wr_ptr_gray[2]~q ),
	.in_wr_ptr_gray_3(\in_wr_ptr_gray[3]~q ),
	.in_wr_ptr_gray_4(\in_wr_ptr_gray[4]~q ),
	.in_wr_ptr_gray_5(\in_wr_ptr_gray[5]~q ),
	.in_wr_ptr_gray_0(\in_wr_ptr_gray[0]~q ));

dffeas \out_rd_ptr_gray[1] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[1]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[1] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[1] .power_up = "low";

dffeas \out_rd_ptr_gray[2] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[2]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[2] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[2] .power_up = "low";

dffeas \out_rd_ptr_gray[3] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[3]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[3] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[3] .power_up = "low";

dffeas \out_rd_ptr_gray[4] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[4]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[4] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[4] .power_up = "low";

dffeas \out_rd_ptr_gray[5] (
	.clk(wire_pll7_clk_1),
	.d(\out_rd_ptr[5]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[5]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[5] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[5] .power_up = "low";

dffeas \out_rd_ptr_gray[0] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[0]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[0] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[0] .power_up = "low";

dffeas \in_wr_ptr_gray[1] (
	.clk(clk_clk),
	.d(\bin2gray~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[1]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[1] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[1] .power_up = "low";

dffeas \in_wr_ptr_gray[2] (
	.clk(clk_clk),
	.d(\bin2gray~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[2]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[2] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[2] .power_up = "low";

dffeas \in_wr_ptr_gray[3] (
	.clk(clk_clk),
	.d(\bin2gray~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[3]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[3] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[3] .power_up = "low";

dffeas \in_wr_ptr_gray[4] (
	.clk(clk_clk),
	.d(\bin2gray~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[4]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[4] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[4] .power_up = "low";

dffeas \in_wr_ptr_gray[5] (
	.clk(clk_clk),
	.d(\in_wr_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[5]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[5] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[5] .power_up = "low";

dffeas \in_wr_ptr_gray[0] (
	.clk(clk_clk),
	.d(\bin2gray~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[0]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[0] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[0] .power_up = "low";

cycloneive_lcell_comb \bin2gray~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[1]~q ),
	.datad(\out_rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\bin2gray~0_combout ),
	.cout());
defparam \bin2gray~0 .lut_mask = 16'h0FF0;
defparam \bin2gray~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[2]~q ),
	.datad(\out_rd_ptr[3]~q ),
	.cin(gnd),
	.combout(\bin2gray~1_combout ),
	.cout());
defparam \bin2gray~1 .lut_mask = 16'h0FF0;
defparam \bin2gray~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[3]~q ),
	.datad(\out_rd_ptr[4]~q ),
	.cin(gnd),
	.combout(\bin2gray~2_combout ),
	.cout());
defparam \bin2gray~2 .lut_mask = 16'h0FF0;
defparam \bin2gray~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[4]~q ),
	.datad(\out_rd_ptr[5]~q ),
	.cin(gnd),
	.combout(\bin2gray~3_combout ),
	.cout());
defparam \bin2gray~3 .lut_mask = 16'h0FF0;
defparam \bin2gray~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[0]~q ),
	.datad(\out_rd_ptr[1]~q ),
	.cin(gnd),
	.combout(\bin2gray~4_combout ),
	.cout());
defparam \bin2gray~4 .lut_mask = 16'h0FF0;
defparam \bin2gray~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[1]~q ),
	.datad(\in_wr_ptr[2]~q ),
	.cin(gnd),
	.combout(\bin2gray~5_combout ),
	.cout());
defparam \bin2gray~5 .lut_mask = 16'h0FF0;
defparam \bin2gray~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[2]~q ),
	.datad(\in_wr_ptr[3]~q ),
	.cin(gnd),
	.combout(\bin2gray~6_combout ),
	.cout());
defparam \bin2gray~6 .lut_mask = 16'h0FF0;
defparam \bin2gray~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[3]~q ),
	.datad(\in_wr_ptr[4]~q ),
	.cin(gnd),
	.combout(\bin2gray~7_combout ),
	.cout());
defparam \bin2gray~7 .lut_mask = 16'h0FF0;
defparam \bin2gray~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[5]~q ),
	.datad(\in_wr_ptr[4]~q ),
	.cin(gnd),
	.combout(\bin2gray~8_combout ),
	.cout());
defparam \bin2gray~8 .lut_mask = 16'h0FF0;
defparam \bin2gray~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[1]~q ),
	.datad(\in_wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\bin2gray~9_combout ),
	.cout());
defparam \bin2gray~9 .lut_mask = 16'h0FF0;
defparam \bin2gray~9 .sum_lutc_input = "datac";

dffeas \out_payload[42] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a18~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_42),
	.prn(vcc));
defparam \out_payload[42] .is_wysiwyg = "true";
defparam \out_payload[42] .power_up = "low";

dffeas \out_payload[43] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a19~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_43),
	.prn(vcc));
defparam \out_payload[43] .is_wysiwyg = "true";
defparam \out_payload[43] .power_up = "low";

dffeas out_valid(
	.clk(wire_pll7_clk_1),
	.d(\empty~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[38] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a17~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_38),
	.prn(vcc));
defparam \out_payload[38] .is_wysiwyg = "true";
defparam \out_payload[38] .power_up = "low";

dffeas \out_payload[37] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a16~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_37),
	.prn(vcc));
defparam \out_payload[37] .is_wysiwyg = "true";
defparam \out_payload[37] .power_up = "low";

dffeas sink_in_reset(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_in_reset1),
	.prn(vcc));
defparam sink_in_reset.is_wysiwyg = "true";
defparam sink_in_reset.power_up = "low";

dffeas full(
	.clk(clk_clk),
	.d(\full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full1),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

dffeas \out_payload[5] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a0~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[6] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a1~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

dffeas \out_payload[7] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a2~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[8] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a3~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

dffeas \out_payload[9] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a4~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_9),
	.prn(vcc));
defparam \out_payload[9] .is_wysiwyg = "true";
defparam \out_payload[9] .power_up = "low";

dffeas \out_payload[10] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a5~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_10),
	.prn(vcc));
defparam \out_payload[10] .is_wysiwyg = "true";
defparam \out_payload[10] .power_up = "low";

dffeas \out_payload[11] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a6~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_11),
	.prn(vcc));
defparam \out_payload[11] .is_wysiwyg = "true";
defparam \out_payload[11] .power_up = "low";

dffeas \out_payload[12] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a7~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[13] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a8~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_13),
	.prn(vcc));
defparam \out_payload[13] .is_wysiwyg = "true";
defparam \out_payload[13] .power_up = "low";

dffeas \out_payload[14] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a9~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_14),
	.prn(vcc));
defparam \out_payload[14] .is_wysiwyg = "true";
defparam \out_payload[14] .power_up = "low";

dffeas \out_payload[15] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a10~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_15),
	.prn(vcc));
defparam \out_payload[15] .is_wysiwyg = "true";
defparam \out_payload[15] .power_up = "low";

dffeas \out_payload[16] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a11~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_16),
	.prn(vcc));
defparam \out_payload[16] .is_wysiwyg = "true";
defparam \out_payload[16] .power_up = "low";

dffeas \out_payload[17] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a12~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_17),
	.prn(vcc));
defparam \out_payload[17] .is_wysiwyg = "true";
defparam \out_payload[17] .power_up = "low";

dffeas \out_payload[18] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a13~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_18),
	.prn(vcc));
defparam \out_payload[18] .is_wysiwyg = "true";
defparam \out_payload[18] .power_up = "low";

dffeas \out_payload[19] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a14~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_19),
	.prn(vcc));
defparam \out_payload[19] .is_wysiwyg = "true";
defparam \out_payload[19] .power_up = "low";

dffeas \out_payload[20] (
	.clk(wire_pll7_clk_1),
	.d(\mem_rtl_0|auto_generated|ram_block1a15~portbdataout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~1_combout ),
	.q(out_payload_20),
	.prn(vcc));
defparam \out_payload[20] .is_wysiwyg = "true";
defparam \out_payload[20] .power_up = "low";

cycloneive_lcell_comb \next_in_wr_ptr~0 (
	.dataa(sink_in_reset1),
	.datab(m0_write),
	.datac(s0_cmd_valid),
	.datad(full1),
	.cin(gnd),
	.combout(\next_in_wr_ptr~0_combout ),
	.cout());
defparam \next_in_wr_ptr~0 .lut_mask = 16'hFEFF;
defparam \next_in_wr_ptr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\in_wr_ptr[0]~q ),
	.datab(\next_in_wr_ptr~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h66EE;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \in_wr_ptr[0] (
	.clk(clk_clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[0]~q ),
	.prn(vcc));
defparam \in_wr_ptr[0] .is_wysiwyg = "true";
defparam \in_wr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\in_wr_ptr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[1] (
	.clk(clk_clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[1]~q ),
	.prn(vcc));
defparam \in_wr_ptr[1] .is_wysiwyg = "true";
defparam \in_wr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \Add0~4 (
	.dataa(\in_wr_ptr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[2] (
	.clk(clk_clk),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[2]~q ),
	.prn(vcc));
defparam \in_wr_ptr[2] .is_wysiwyg = "true";
defparam \in_wr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add0~6 (
	.dataa(\in_wr_ptr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[3] (
	.clk(clk_clk),
	.d(\Add0~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[3]~q ),
	.prn(vcc));
defparam \in_wr_ptr[3] .is_wysiwyg = "true";
defparam \in_wr_ptr[3] .power_up = "low";

cycloneive_lcell_comb \Add0~8 (
	.dataa(\in_wr_ptr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[4] (
	.clk(clk_clk),
	.d(\Add0~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[4]~q ),
	.prn(vcc));
defparam \in_wr_ptr[4] .is_wysiwyg = "true";
defparam \in_wr_ptr[4] .power_up = "low";

dffeas \out_rd_ptr[0] (
	.clk(wire_pll7_clk_1),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[0]~q ),
	.prn(vcc));
defparam \out_rd_ptr[0] .is_wysiwyg = "true";
defparam \out_rd_ptr[0] .power_up = "low";

cycloneive_lcell_comb \internal_out_ready~0 (
	.dataa(old_read),
	.datab(gnd),
	.datac(stop_cmd_r),
	.datad(out_payload_38),
	.cin(gnd),
	.combout(\internal_out_ready~0_combout ),
	.cout());
defparam \internal_out_ready~0 .lut_mask = 16'hAFFF;
defparam \internal_out_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_ready~1 (
	.dataa(\internal_out_ready~0_combout ),
	.datab(waitrequest_reset_override),
	.datac(av_waitrequest_generated),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_ready~1_combout ),
	.cout());
defparam \internal_out_ready~1 .lut_mask = 16'hEFFF;
defparam \internal_out_ready~1 .sum_lutc_input = "datac";

dffeas \out_rd_ptr[1] (
	.clk(wire_pll7_clk_1),
	.d(\Add1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[1]~q ),
	.prn(vcc));
defparam \out_rd_ptr[1] .is_wysiwyg = "true";
defparam \out_rd_ptr[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\out_rd_ptr[0]~q ),
	.datab(\next_out_rd_ptr~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
defparam \Add1~0 .lut_mask = 16'h66EE;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~2 (
	.dataa(\out_rd_ptr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\write_crosser|sync[4].u|dreg[1]~q ),
	.datad(\write_crosser|sync[5].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h0FF0;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\write_crosser|sync[1].u|dreg[1]~q ),
	.datab(\write_crosser|sync[2].u|dreg[1]~q ),
	.datac(\write_crosser|sync[3].u|dreg[1]~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\Add1~2_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Add1~0_combout ),
	.datad(\write_crosser|sync[0].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h6996;
defparam \Equal0~2 .sum_lutc_input = "datac";

dffeas \out_rd_ptr[4] (
	.clk(wire_pll7_clk_1),
	.d(\Add1~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[4]~q ),
	.prn(vcc));
defparam \out_rd_ptr[4] .is_wysiwyg = "true";
defparam \out_rd_ptr[4] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(\out_rd_ptr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
defparam \Add1~4 .lut_mask = 16'h5AAF;
defparam \Add1~4 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[2] (
	.clk(wire_pll7_clk_1),
	.d(\Add1~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[2]~q ),
	.prn(vcc));
defparam \out_rd_ptr[2] .is_wysiwyg = "true";
defparam \out_rd_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(\out_rd_ptr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[3] (
	.clk(wire_pll7_clk_1),
	.d(\Add1~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[3]~q ),
	.prn(vcc));
defparam \out_rd_ptr[3] .is_wysiwyg = "true";
defparam \out_rd_ptr[3] .power_up = "low";

cycloneive_lcell_comb \Add1~8 (
	.dataa(\out_rd_ptr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
defparam \Add1~8 .lut_mask = 16'h5AAF;
defparam \Add1~8 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[5] (
	.clk(wire_pll7_clk_1),
	.d(\Add1~10_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[5]~q ),
	.prn(vcc));
defparam \out_rd_ptr[5] .is_wysiwyg = "true";
defparam \out_rd_ptr[5] .power_up = "low";

cycloneive_lcell_comb \Add1~10 (
	.dataa(\out_rd_ptr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\write_crosser|sync[4].u|dreg[1]~q ),
	.datab(\write_crosser|sync[5].u|dreg[1]~q ),
	.datac(\Add1~8_combout ),
	.datad(\Add1~10_combout ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h6996;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\Add1~4_combout ),
	.datab(\write_crosser|sync[2].u|dreg[1]~q ),
	.datac(\write_crosser|sync[3].u|dreg[1]~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'h6996;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\write_crosser|sync[4].u|dreg[1]~q ),
	.datab(\write_crosser|sync[5].u|dreg[1]~q ),
	.datac(\Add1~6_combout ),
	.datad(\write_crosser|sync[3].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'h6996;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\Equal0~4_combout ),
	.datad(\Equal0~5_combout ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hFFF7;
defparam \Equal0~6 .sum_lutc_input = "datac";

dffeas empty(
	.clk(wire_pll7_clk_1),
	.d(\Equal0~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

cycloneive_lcell_comb \next_out_rd_ptr~0 (
	.dataa(\internal_out_ready~1_combout ),
	.datab(\empty~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_out_rd_ptr~0_combout ),
	.cout());
defparam \next_out_rd_ptr~0 .lut_mask = 16'hEEEE;
defparam \next_out_rd_ptr~0 .sum_lutc_input = "datac";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a18 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,W_alu_result_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a18 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_first_bit_number = 18;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_first_bit_number = 18;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a19 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,W_alu_result_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a19 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_first_bit_number = 19;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_first_bit_number = 19;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a17 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,m0_read}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a17 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_first_bit_number = 17;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_first_bit_number = 17;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a16 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,m0_write1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a16 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_first_bit_number = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_first_bit_number = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .ram_block_type = "auto";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\read_crosser|sync[4].u|dreg[1]~q ),
	.datad(\read_crosser|sync[5].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h0FF0;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(\read_crosser|sync[1].u|dreg[1]~q ),
	.datab(\read_crosser|sync[2].u|dreg[1]~q ),
	.datac(\read_crosser|sync[3].u|dreg[1]~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h6996;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~0 (
	.dataa(\Add0~2_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Add0~0_combout ),
	.datad(\read_crosser|sync[0].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\full~0_combout ),
	.cout());
defparam \full~0 .lut_mask = 16'h6996;
defparam \full~0 .sum_lutc_input = "datac";

dffeas \in_wr_ptr[5] (
	.clk(clk_clk),
	.d(\Add0~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[5]~q ),
	.prn(vcc));
defparam \in_wr_ptr[5] .is_wysiwyg = "true";
defparam \in_wr_ptr[5] .power_up = "low";

cycloneive_lcell_comb \Add0~10 (
	.dataa(\in_wr_ptr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout());
defparam \Add0~10 .lut_mask = 16'h5A5A;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \full~1 (
	.dataa(\read_crosser|sync[4].u|dreg[1]~q ),
	.datab(\read_crosser|sync[5].u|dreg[1]~q ),
	.datac(\Add0~8_combout ),
	.datad(\Add0~10_combout ),
	.cin(gnd),
	.combout(\full~1_combout ),
	.cout());
defparam \full~1 .lut_mask = 16'h6996;
defparam \full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(\read_crosser|sync[2].u|dreg[1]~q ),
	.datab(\read_crosser|sync[3].u|dreg[1]~q ),
	.datac(\Equal1~0_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'h6996;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~3 (
	.dataa(\read_crosser|sync[4].u|dreg[1]~q ),
	.datab(\read_crosser|sync[5].u|dreg[1]~q ),
	.datac(\read_crosser|sync[3].u|dreg[1]~q ),
	.datad(\Add0~6_combout ),
	.cin(gnd),
	.combout(\Equal1~3_combout ),
	.cout());
defparam \Equal1~3 .lut_mask = 16'h6996;
defparam \Equal1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~2 (
	.dataa(\full~0_combout ),
	.datab(\full~1_combout ),
	.datac(\Equal1~2_combout ),
	.datad(\Equal1~3_combout ),
	.cin(gnd),
	.combout(\full~2_combout ),
	.cout());
defparam \full~2 .lut_mask = 16'hEFFF;
defparam \full~2 .sum_lutc_input = "datac";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a0 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a1 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a2 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a3 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a4 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a5 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a6 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a7 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a8 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_8}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a8 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_first_bit_number = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_first_bit_number = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a9 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_9}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a9 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_first_bit_number = 9;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_first_bit_number = 9;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a10 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_10}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a10 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_first_bit_number = 10;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_first_bit_number = 10;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a11 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a11 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_first_bit_number = 11;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_first_bit_number = 11;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a12 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_12}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a12 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_first_bit_number = 12;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_first_bit_number = 12;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a13 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_13}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a13 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_first_bit_number = 13;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_first_bit_number = 13;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a14 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_14}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a14 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_first_bit_number = 14;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_first_bit_number = 14;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a15 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk_clk),
	.clk1(wire_pll7_clk_1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_15}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a15 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:cmd_fifo|altsyncram:mem_rtl_0|altsyncram_evc1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_first_bit_number = 15;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_width = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_first_bit_number = 15;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_last_address = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_depth = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_width = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .ram_block_type = "auto";

endmodule

module usb_system_altera_dcfifo_synchronizer_bundle (
	r_sync_rst,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	out_rd_ptr_gray_1,
	out_rd_ptr_gray_2,
	out_rd_ptr_gray_3,
	out_rd_ptr_gray_4,
	out_rd_ptr_gray_5,
	out_rd_ptr_gray_0,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
input 	out_rd_ptr_gray_1;
input 	out_rd_ptr_gray_2;
input 	out_rd_ptr_gray_3;
input 	out_rd_ptr_gray_4;
input 	out_rd_ptr_gray_5;
input 	out_rd_ptr_gray_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_std_synchronizer_nocut_5 \sync[5].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_14),
	.din(out_rd_ptr_gray_5),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_4 \sync[4].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_13),
	.din(out_rd_ptr_gray_4),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_3 \sync[3].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_12),
	.din(out_rd_ptr_gray_3),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_2 \sync[2].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_11),
	.din(out_rd_ptr_gray_2),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_1 \sync[1].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_1),
	.din(out_rd_ptr_gray_1),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut \sync[0].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_15),
	.din(out_rd_ptr_gray_0),
	.clk(clk_clk));

endmodule

module usb_system_altera_std_synchronizer_nocut (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_1 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_2 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_3 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_4 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_5 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_dcfifo_synchronizer_bundle_1 (
	wire_pll7_clk_1,
	altera_reset_synchronizer_int_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	in_wr_ptr_gray_1,
	in_wr_ptr_gray_2,
	in_wr_ptr_gray_3,
	in_wr_ptr_gray_4,
	in_wr_ptr_gray_5,
	in_wr_ptr_gray_0)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
input 	altera_reset_synchronizer_int_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
input 	in_wr_ptr_gray_1;
input 	in_wr_ptr_gray_2;
input 	in_wr_ptr_gray_3;
input 	in_wr_ptr_gray_4;
input 	in_wr_ptr_gray_5;
input 	in_wr_ptr_gray_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_std_synchronizer_nocut_11 \sync[5].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_14),
	.din(in_wr_ptr_gray_5));

usb_system_altera_std_synchronizer_nocut_10 \sync[4].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_13),
	.din(in_wr_ptr_gray_4));

usb_system_altera_std_synchronizer_nocut_9 \sync[3].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_12),
	.din(in_wr_ptr_gray_3));

usb_system_altera_std_synchronizer_nocut_8 \sync[2].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_11),
	.din(in_wr_ptr_gray_2));

usb_system_altera_std_synchronizer_nocut_7 \sync[1].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_1),
	.din(in_wr_ptr_gray_1));

usb_system_altera_std_synchronizer_nocut_6 \sync[0].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_15),
	.din(in_wr_ptr_gray_0));

endmodule

module usb_system_altera_std_synchronizer_nocut_6 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_7 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_8 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_9 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_10 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_11 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_avalon_dc_fifo_1 (
	wire_pll7_clk_1,
	in_space_avail_8,
	in_space_avail_7,
	in_space_avail_6,
	in_space_avail_5,
	in_space_avail_4,
	in_space_avail_3,
	in_space_avail_2,
	in_space_avail_1,
	in_space_avail_0,
	altera_reset_synchronizer_int_chain_out,
	r_sync_rst,
	out_valid1,
	read_latency_shift_reg_0,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_5,
	out_payload_6,
	out_payload_7,
	out_payload_8,
	out_payload_9,
	out_payload_10,
	out_payload_11,
	out_payload_12,
	out_payload_13,
	out_payload_14,
	out_payload_15,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
output 	in_space_avail_8;
output 	in_space_avail_7;
output 	in_space_avail_6;
output 	in_space_avail_5;
output 	in_space_avail_4;
output 	in_space_avail_3;
output 	in_space_avail_2;
output 	in_space_avail_1;
output 	in_space_avail_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	r_sync_rst;
output 	out_valid1;
input 	read_latency_shift_reg_0;
output 	out_payload_0;
output 	out_payload_1;
output 	out_payload_2;
output 	out_payload_3;
output 	out_payload_4;
output 	out_payload_5;
output 	out_payload_6;
output 	out_payload_7;
output 	out_payload_8;
output 	out_payload_9;
output 	out_payload_10;
output 	out_payload_11;
output 	out_payload_12;
output 	out_payload_13;
output 	out_payload_14;
output 	out_payload_15;
input 	av_readdata_pre_0;
input 	av_readdata_pre_1;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_6;
input 	av_readdata_pre_7;
input 	av_readdata_pre_8;
input 	av_readdata_pre_9;
input 	av_readdata_pre_10;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_crosser|sync[8].u|dreg[1]~q ;
wire \read_crosser|sync[7].u|dreg[1]~q ;
wire \read_crosser|sync[6].u|dreg[1]~q ;
wire \read_crosser|sync[5].u|dreg[1]~q ;
wire \read_crosser|sync[4].u|dreg[1]~q ;
wire \read_crosser|sync[3].u|dreg[1]~q ;
wire \read_crosser|sync[2].u|dreg[1]~q ;
wire \read_crosser|sync[1].u|dreg[1]~q ;
wire \read_crosser|sync[0].u|dreg[1]~q ;
wire \write_crosser|sync[0].u|dreg[1]~q ;
wire \write_crosser|sync[1].u|dreg[1]~q ;
wire \write_crosser|sync[2].u|dreg[1]~q ;
wire \write_crosser|sync[3].u|dreg[1]~q ;
wire \write_crosser|sync[4].u|dreg[1]~q ;
wire \write_crosser|sync[5].u|dreg[1]~q ;
wire \write_crosser|sync[6].u|dreg[1]~q ;
wire \write_crosser|sync[7].u|dreg[1]~q ;
wire \write_crosser|sync[8].u|dreg[1]~q ;
wire \out_rd_ptr_gray[8]~q ;
wire \out_rd_ptr_gray[7]~q ;
wire \out_rd_ptr_gray[6]~q ;
wire \out_rd_ptr_gray[5]~q ;
wire \out_rd_ptr_gray[4]~q ;
wire \out_rd_ptr_gray[3]~q ;
wire \out_rd_ptr_gray[2]~q ;
wire \out_rd_ptr_gray[1]~q ;
wire \out_rd_ptr_gray[0]~q ;
wire \in_wr_ptr_gray[0]~q ;
wire \in_wr_ptr_gray[1]~q ;
wire \in_wr_ptr_gray[2]~q ;
wire \in_wr_ptr_gray[3]~q ;
wire \in_wr_ptr_gray[4]~q ;
wire \in_wr_ptr_gray[5]~q ;
wire \in_wr_ptr_gray[6]~q ;
wire \in_wr_ptr_gray[7]~q ;
wire \in_wr_ptr_gray[8]~q ;
wire \bin2gray~0_combout ;
wire \bin2gray~1_combout ;
wire \bin2gray~2_combout ;
wire \bin2gray~3_combout ;
wire \bin2gray~4_combout ;
wire \bin2gray~5_combout ;
wire \bin2gray~6_combout ;
wire \bin2gray~7_combout ;
wire \bin2gray~8_combout ;
wire \bin2gray~9_combout ;
wire \bin2gray~10_combout ;
wire \bin2gray~11_combout ;
wire \bin2gray~12_combout ;
wire \bin2gray~13_combout ;
wire \bin2gray~14_combout ;
wire \bin2gray~15_combout ;
wire \in_wr_ptr[8]~q ;
wire \next_in_rd_ptr[5]~2_combout ;
wire \next_in_rd_ptr[1]~5_combout ;
wire \full~0_combout ;
wire \full~1_combout ;
wire \full~2_combout ;
wire \next_in_rd_ptr[5]~1_combout ;
wire \full~3_combout ;
wire \next_in_rd_ptr[3]~4_combout ;
wire \full~4_combout ;
wire \next_in_rd_ptr[0]~combout ;
wire \full~5_combout ;
wire \full~q ;
wire \next_in_wr_ptr~0_combout ;
wire \Add0~0_combout ;
wire \in_wr_ptr[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \in_wr_ptr[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \in_wr_ptr[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \in_wr_ptr[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \in_wr_ptr[4]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \in_wr_ptr[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \in_wr_ptr[6]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \in_wr_ptr[7]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \next_in_rd_ptr[7]~0_combout ;
wire \next_in_rd_ptr[3]~3_combout ;
wire \next_in_rd_ptr[0]~6_combout ;
wire \in_space_avail[0]~10 ;
wire \in_space_avail[1]~12 ;
wire \in_space_avail[2]~14 ;
wire \in_space_avail[3]~16 ;
wire \in_space_avail[4]~18 ;
wire \in_space_avail[5]~20 ;
wire \in_space_avail[6]~22 ;
wire \in_space_avail[7]~24 ;
wire \in_space_avail[8]~25_combout ;
wire \in_space_avail[7]~23_combout ;
wire \in_space_avail[6]~21_combout ;
wire \in_space_avail[5]~19_combout ;
wire \in_space_avail[4]~17_combout ;
wire \in_space_avail[3]~15_combout ;
wire \in_space_avail[2]~13_combout ;
wire \in_space_avail[1]~11_combout ;
wire \in_space_avail[0]~9_combout ;
wire \out_rd_ptr[1]~q ;
wire \Add1~0_combout ;
wire \out_rd_ptr[0]~q ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \out_rd_ptr[8]~q ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \out_rd_ptr[2]~q ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \out_rd_ptr[3]~q ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \out_rd_ptr[4]~q ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \out_rd_ptr[5]~q ;
wire \Add1~11 ;
wire \Add1~12_combout ;
wire \out_rd_ptr[6]~q ;
wire \Add1~13 ;
wire \Add1~14_combout ;
wire \out_rd_ptr[7]~q ;
wire \Add1~15 ;
wire \Add1~16_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Equal0~6_combout ;
wire \Equal0~7_combout ;
wire \Equal0~8_combout ;
wire \Equal0~9_combout ;
wire \empty~q ;
wire \mem_rtl_0|auto_generated|ram_block1a0~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a1~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a2~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a3~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a4~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a5~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a6~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a7~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a8~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a9~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a10~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a11~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a12~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a13~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a14~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a15~portbdataout ;

wire [143:0] \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ;

assign \mem_rtl_0|auto_generated|ram_block1a0~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a1~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a2~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a3~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a4~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a5~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a6~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a7~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a8~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a9~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a10~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a11~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a12~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a13~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a14~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a15~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus [0];

usb_system_altera_dcfifo_synchronizer_bundle_2 read_crosser(
	.wire_pll7_clk_1(wire_pll7_clk_1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.dreg_1(\read_crosser|sync[8].u|dreg[1]~q ),
	.dreg_11(\read_crosser|sync[7].u|dreg[1]~q ),
	.dreg_12(\read_crosser|sync[6].u|dreg[1]~q ),
	.dreg_13(\read_crosser|sync[5].u|dreg[1]~q ),
	.dreg_14(\read_crosser|sync[4].u|dreg[1]~q ),
	.dreg_15(\read_crosser|sync[3].u|dreg[1]~q ),
	.dreg_16(\read_crosser|sync[2].u|dreg[1]~q ),
	.dreg_17(\read_crosser|sync[1].u|dreg[1]~q ),
	.dreg_18(\read_crosser|sync[0].u|dreg[1]~q ),
	.out_rd_ptr_gray_8(\out_rd_ptr_gray[8]~q ),
	.out_rd_ptr_gray_7(\out_rd_ptr_gray[7]~q ),
	.out_rd_ptr_gray_6(\out_rd_ptr_gray[6]~q ),
	.out_rd_ptr_gray_5(\out_rd_ptr_gray[5]~q ),
	.out_rd_ptr_gray_4(\out_rd_ptr_gray[4]~q ),
	.out_rd_ptr_gray_3(\out_rd_ptr_gray[3]~q ),
	.out_rd_ptr_gray_2(\out_rd_ptr_gray[2]~q ),
	.out_rd_ptr_gray_1(\out_rd_ptr_gray[1]~q ),
	.out_rd_ptr_gray_0(\out_rd_ptr_gray[0]~q ));

usb_system_altera_dcfifo_synchronizer_bundle_3 write_crosser(
	.r_sync_rst(r_sync_rst),
	.dreg_1(\write_crosser|sync[0].u|dreg[1]~q ),
	.dreg_11(\write_crosser|sync[1].u|dreg[1]~q ),
	.dreg_12(\write_crosser|sync[2].u|dreg[1]~q ),
	.dreg_13(\write_crosser|sync[3].u|dreg[1]~q ),
	.dreg_14(\write_crosser|sync[4].u|dreg[1]~q ),
	.dreg_15(\write_crosser|sync[5].u|dreg[1]~q ),
	.dreg_16(\write_crosser|sync[6].u|dreg[1]~q ),
	.dreg_17(\write_crosser|sync[7].u|dreg[1]~q ),
	.dreg_18(\write_crosser|sync[8].u|dreg[1]~q ),
	.in_wr_ptr_gray_0(\in_wr_ptr_gray[0]~q ),
	.in_wr_ptr_gray_1(\in_wr_ptr_gray[1]~q ),
	.in_wr_ptr_gray_2(\in_wr_ptr_gray[2]~q ),
	.in_wr_ptr_gray_3(\in_wr_ptr_gray[3]~q ),
	.in_wr_ptr_gray_4(\in_wr_ptr_gray[4]~q ),
	.in_wr_ptr_gray_5(\in_wr_ptr_gray[5]~q ),
	.in_wr_ptr_gray_6(\in_wr_ptr_gray[6]~q ),
	.in_wr_ptr_gray_7(\in_wr_ptr_gray[7]~q ),
	.in_wr_ptr_gray_8(\in_wr_ptr_gray[8]~q ),
	.clk_clk(clk_clk));

dffeas \out_rd_ptr_gray[8] (
	.clk(clk_clk),
	.d(\out_rd_ptr[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[8]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[8] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[8] .power_up = "low";

dffeas \out_rd_ptr_gray[7] (
	.clk(clk_clk),
	.d(\bin2gray~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[7]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[7] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[7] .power_up = "low";

dffeas \out_rd_ptr_gray[6] (
	.clk(clk_clk),
	.d(\bin2gray~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[6]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[6] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[6] .power_up = "low";

dffeas \out_rd_ptr_gray[5] (
	.clk(clk_clk),
	.d(\bin2gray~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[5]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[5] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[5] .power_up = "low";

dffeas \out_rd_ptr_gray[4] (
	.clk(clk_clk),
	.d(\bin2gray~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[4]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[4] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[4] .power_up = "low";

dffeas \out_rd_ptr_gray[3] (
	.clk(clk_clk),
	.d(\bin2gray~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[3]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[3] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[3] .power_up = "low";

dffeas \out_rd_ptr_gray[2] (
	.clk(clk_clk),
	.d(\bin2gray~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[2]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[2] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[2] .power_up = "low";

dffeas \out_rd_ptr_gray[1] (
	.clk(clk_clk),
	.d(\bin2gray~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[1]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[1] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[1] .power_up = "low";

dffeas \out_rd_ptr_gray[0] (
	.clk(clk_clk),
	.d(\bin2gray~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr_gray[0]~q ),
	.prn(vcc));
defparam \out_rd_ptr_gray[0] .is_wysiwyg = "true";
defparam \out_rd_ptr_gray[0] .power_up = "low";

dffeas \in_wr_ptr_gray[0] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[0]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[0] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[0] .power_up = "low";

dffeas \in_wr_ptr_gray[1] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[1]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[1] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[1] .power_up = "low";

dffeas \in_wr_ptr_gray[2] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~10_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[2]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[2] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[2] .power_up = "low";

dffeas \in_wr_ptr_gray[3] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~11_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[3]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[3] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[3] .power_up = "low";

dffeas \in_wr_ptr_gray[4] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[4]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[4] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[4] .power_up = "low";

dffeas \in_wr_ptr_gray[5] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[5]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[5] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[5] .power_up = "low";

dffeas \in_wr_ptr_gray[6] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~14_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[6]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[6] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[6] .power_up = "low";

dffeas \in_wr_ptr_gray[7] (
	.clk(wire_pll7_clk_1),
	.d(\bin2gray~15_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[7]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[7] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[7] .power_up = "low";

dffeas \in_wr_ptr_gray[8] (
	.clk(wire_pll7_clk_1),
	.d(\in_wr_ptr[8]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr_gray[8]~q ),
	.prn(vcc));
defparam \in_wr_ptr_gray[8] .is_wysiwyg = "true";
defparam \in_wr_ptr_gray[8] .power_up = "low";

cycloneive_lcell_comb \bin2gray~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[7]~q ),
	.datad(\out_rd_ptr[8]~q ),
	.cin(gnd),
	.combout(\bin2gray~0_combout ),
	.cout());
defparam \bin2gray~0 .lut_mask = 16'h0FF0;
defparam \bin2gray~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[6]~q ),
	.datad(\out_rd_ptr[7]~q ),
	.cin(gnd),
	.combout(\bin2gray~1_combout ),
	.cout());
defparam \bin2gray~1 .lut_mask = 16'h0FF0;
defparam \bin2gray~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[6]~q ),
	.datad(\out_rd_ptr[5]~q ),
	.cin(gnd),
	.combout(\bin2gray~2_combout ),
	.cout());
defparam \bin2gray~2 .lut_mask = 16'h0FF0;
defparam \bin2gray~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[5]~q ),
	.datad(\out_rd_ptr[4]~q ),
	.cin(gnd),
	.combout(\bin2gray~3_combout ),
	.cout());
defparam \bin2gray~3 .lut_mask = 16'h0FF0;
defparam \bin2gray~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[4]~q ),
	.datad(\out_rd_ptr[3]~q ),
	.cin(gnd),
	.combout(\bin2gray~4_combout ),
	.cout());
defparam \bin2gray~4 .lut_mask = 16'h0FF0;
defparam \bin2gray~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[3]~q ),
	.datad(\out_rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\bin2gray~5_combout ),
	.cout());
defparam \bin2gray~5 .lut_mask = 16'h0FF0;
defparam \bin2gray~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[1]~q ),
	.datad(\out_rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\bin2gray~6_combout ),
	.cout());
defparam \bin2gray~6 .lut_mask = 16'h0FF0;
defparam \bin2gray~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_rd_ptr[1]~q ),
	.datad(\out_rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\bin2gray~7_combout ),
	.cout());
defparam \bin2gray~7 .lut_mask = 16'h0FF0;
defparam \bin2gray~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[1]~q ),
	.datad(\in_wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\bin2gray~8_combout ),
	.cout());
defparam \bin2gray~8 .lut_mask = 16'h0FF0;
defparam \bin2gray~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[2]~q ),
	.datad(\in_wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\bin2gray~9_combout ),
	.cout());
defparam \bin2gray~9 .lut_mask = 16'h0FF0;
defparam \bin2gray~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[3]~q ),
	.datad(\in_wr_ptr[2]~q ),
	.cin(gnd),
	.combout(\bin2gray~10_combout ),
	.cout());
defparam \bin2gray~10 .lut_mask = 16'h0FF0;
defparam \bin2gray~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[4]~q ),
	.datad(\in_wr_ptr[3]~q ),
	.cin(gnd),
	.combout(\bin2gray~11_combout ),
	.cout());
defparam \bin2gray~11 .lut_mask = 16'h0FF0;
defparam \bin2gray~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[5]~q ),
	.datad(\in_wr_ptr[4]~q ),
	.cin(gnd),
	.combout(\bin2gray~12_combout ),
	.cout());
defparam \bin2gray~12 .lut_mask = 16'h0FF0;
defparam \bin2gray~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[6]~q ),
	.datad(\in_wr_ptr[5]~q ),
	.cin(gnd),
	.combout(\bin2gray~13_combout ),
	.cout());
defparam \bin2gray~13 .lut_mask = 16'h0FF0;
defparam \bin2gray~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[7]~q ),
	.datad(\in_wr_ptr[6]~q ),
	.cin(gnd),
	.combout(\bin2gray~14_combout ),
	.cout());
defparam \bin2gray~14 .lut_mask = 16'h0FF0;
defparam \bin2gray~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bin2gray~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_wr_ptr[8]~q ),
	.datad(\in_wr_ptr[7]~q ),
	.cin(gnd),
	.combout(\bin2gray~15_combout ),
	.cout());
defparam \bin2gray~15 .lut_mask = 16'h0FF0;
defparam \bin2gray~15 .sum_lutc_input = "datac";

dffeas \in_space_avail[8] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[8]~25_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_8),
	.prn(vcc));
defparam \in_space_avail[8] .is_wysiwyg = "true";
defparam \in_space_avail[8] .power_up = "low";

dffeas \in_space_avail[7] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[7]~23_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_7),
	.prn(vcc));
defparam \in_space_avail[7] .is_wysiwyg = "true";
defparam \in_space_avail[7] .power_up = "low";

dffeas \in_space_avail[6] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[6]~21_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_6),
	.prn(vcc));
defparam \in_space_avail[6] .is_wysiwyg = "true";
defparam \in_space_avail[6] .power_up = "low";

dffeas \in_space_avail[5] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[5]~19_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_5),
	.prn(vcc));
defparam \in_space_avail[5] .is_wysiwyg = "true";
defparam \in_space_avail[5] .power_up = "low";

dffeas \in_space_avail[4] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[4]~17_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_4),
	.prn(vcc));
defparam \in_space_avail[4] .is_wysiwyg = "true";
defparam \in_space_avail[4] .power_up = "low";

dffeas \in_space_avail[3] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[3]~15_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_3),
	.prn(vcc));
defparam \in_space_avail[3] .is_wysiwyg = "true";
defparam \in_space_avail[3] .power_up = "low";

dffeas \in_space_avail[2] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[2]~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_2),
	.prn(vcc));
defparam \in_space_avail[2] .is_wysiwyg = "true";
defparam \in_space_avail[2] .power_up = "low";

dffeas \in_space_avail[1] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[1]~11_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_1),
	.prn(vcc));
defparam \in_space_avail[1] .is_wysiwyg = "true";
defparam \in_space_avail[1] .power_up = "low";

dffeas \in_space_avail[0] (
	.clk(wire_pll7_clk_1),
	.d(\in_space_avail[0]~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_space_avail_0),
	.prn(vcc));
defparam \in_space_avail[0] .is_wysiwyg = "true";
defparam \in_space_avail[0] .power_up = "low";

dffeas out_valid(
	.clk(clk_clk),
	.d(\empty~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[0] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a0~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a1~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a2~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas \out_payload[3] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a3~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_3),
	.prn(vcc));
defparam \out_payload[3] .is_wysiwyg = "true";
defparam \out_payload[3] .power_up = "low";

dffeas \out_payload[4] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a4~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_4),
	.prn(vcc));
defparam \out_payload[4] .is_wysiwyg = "true";
defparam \out_payload[4] .power_up = "low";

dffeas \out_payload[5] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a5~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[6] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a6~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

dffeas \out_payload[7] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a7~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[8] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a8~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

dffeas \out_payload[9] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a9~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_9),
	.prn(vcc));
defparam \out_payload[9] .is_wysiwyg = "true";
defparam \out_payload[9] .power_up = "low";

dffeas \out_payload[10] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a10~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_10),
	.prn(vcc));
defparam \out_payload[10] .is_wysiwyg = "true";
defparam \out_payload[10] .power_up = "low";

dffeas \out_payload[11] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a11~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_11),
	.prn(vcc));
defparam \out_payload[11] .is_wysiwyg = "true";
defparam \out_payload[11] .power_up = "low";

dffeas \out_payload[12] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a12~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[13] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a13~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_13),
	.prn(vcc));
defparam \out_payload[13] .is_wysiwyg = "true";
defparam \out_payload[13] .power_up = "low";

dffeas \out_payload[14] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a14~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_14),
	.prn(vcc));
defparam \out_payload[14] .is_wysiwyg = "true";
defparam \out_payload[14] .power_up = "low";

dffeas \out_payload[15] (
	.clk(clk_clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a15~portbdataout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_payload_15),
	.prn(vcc));
defparam \out_payload[15] .is_wysiwyg = "true";
defparam \out_payload[15] .power_up = "low";

dffeas \in_wr_ptr[8] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~16_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[8]~q ),
	.prn(vcc));
defparam \in_wr_ptr[8] .is_wysiwyg = "true";
defparam \in_wr_ptr[8] .power_up = "low";

cycloneive_lcell_comb \next_in_rd_ptr[5]~2 (
	.dataa(\read_crosser|sync[8].u|dreg[1]~q ),
	.datab(\read_crosser|sync[7].u|dreg[1]~q ),
	.datac(\read_crosser|sync[6].u|dreg[1]~q ),
	.datad(\read_crosser|sync[5].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\next_in_rd_ptr[5]~2_combout ),
	.cout());
defparam \next_in_rd_ptr[5]~2 .lut_mask = 16'h6996;
defparam \next_in_rd_ptr[5]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_in_rd_ptr[1]~5 (
	.dataa(\next_in_rd_ptr[5]~2_combout ),
	.datab(\read_crosser|sync[4].u|dreg[1]~q ),
	.datac(\read_crosser|sync[3].u|dreg[1]~q ),
	.datad(\read_crosser|sync[2].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\next_in_rd_ptr[1]~5_combout ),
	.cout());
defparam \next_in_rd_ptr[1]~5 .lut_mask = 16'h6996;
defparam \next_in_rd_ptr[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~0 (
	.dataa(\Add0~4_combout ),
	.datab(\next_in_rd_ptr[1]~5_combout ),
	.datac(\Add0~2_combout ),
	.datad(\read_crosser|sync[1].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\full~0_combout ),
	.cout());
defparam \full~0 .lut_mask = 16'h6996;
defparam \full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~1 (
	.dataa(\Add0~10_combout ),
	.datab(\next_in_rd_ptr[5]~2_combout ),
	.datac(\Add0~8_combout ),
	.datad(\read_crosser|sync[4].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\full~1_combout ),
	.cout());
defparam \full~1 .lut_mask = 16'h6996;
defparam \full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~2 (
	.dataa(\Add0~14_combout ),
	.datab(\read_crosser|sync[7].u|dreg[1]~q ),
	.datac(\Add0~16_combout ),
	.datad(\read_crosser|sync[8].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\full~2_combout ),
	.cout());
defparam \full~2 .lut_mask = 16'h6996;
defparam \full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_in_rd_ptr[5]~1 (
	.dataa(\read_crosser|sync[8].u|dreg[1]~q ),
	.datab(\read_crosser|sync[7].u|dreg[1]~q ),
	.datac(\read_crosser|sync[6].u|dreg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_in_rd_ptr[5]~1_combout ),
	.cout());
defparam \next_in_rd_ptr[5]~1 .lut_mask = 16'h9696;
defparam \next_in_rd_ptr[5]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~3 (
	.dataa(\full~1_combout ),
	.datab(\full~2_combout ),
	.datac(\Add0~12_combout ),
	.datad(\next_in_rd_ptr[5]~1_combout ),
	.cin(gnd),
	.combout(\full~3_combout ),
	.cout());
defparam \full~3 .lut_mask = 16'hEFFE;
defparam \full~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_in_rd_ptr[3]~4 (
	.dataa(\next_in_rd_ptr[5]~2_combout ),
	.datab(\read_crosser|sync[4].u|dreg[1]~q ),
	.datac(\read_crosser|sync[3].u|dreg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_in_rd_ptr[3]~4_combout ),
	.cout());
defparam \next_in_rd_ptr[3]~4 .lut_mask = 16'h9696;
defparam \next_in_rd_ptr[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~4 (
	.dataa(\full~0_combout ),
	.datab(\full~3_combout ),
	.datac(\Add0~6_combout ),
	.datad(\next_in_rd_ptr[3]~4_combout ),
	.cin(gnd),
	.combout(\full~4_combout ),
	.cout());
defparam \full~4 .lut_mask = 16'hEFFE;
defparam \full~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_in_rd_ptr[0] (
	.dataa(\next_in_rd_ptr[1]~5_combout ),
	.datab(\read_crosser|sync[1].u|dreg[1]~q ),
	.datac(\read_crosser|sync[0].u|dreg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_in_rd_ptr[0]~combout ),
	.cout());
defparam \next_in_rd_ptr[0] .lut_mask = 16'h9696;
defparam \next_in_rd_ptr[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \full~5 (
	.dataa(\full~4_combout ),
	.datab(\Add0~0_combout ),
	.datac(\next_in_rd_ptr[0]~combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\full~5_combout ),
	.cout());
defparam \full~5 .lut_mask = 16'hBEBE;
defparam \full~5 .sum_lutc_input = "datac";

dffeas full(
	.clk(wire_pll7_clk_1),
	.d(\full~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\full~q ),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

cycloneive_lcell_comb \next_in_wr_ptr~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\full~q ),
	.cin(gnd),
	.combout(\next_in_wr_ptr~0_combout ),
	.cout());
defparam \next_in_wr_ptr~0 .lut_mask = 16'hAAFF;
defparam \next_in_wr_ptr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\in_wr_ptr[0]~q ),
	.datab(\next_in_wr_ptr~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h66EE;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \in_wr_ptr[0] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[0]~q ),
	.prn(vcc));
defparam \in_wr_ptr[0] .is_wysiwyg = "true";
defparam \in_wr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\in_wr_ptr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[1] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[1]~q ),
	.prn(vcc));
defparam \in_wr_ptr[1] .is_wysiwyg = "true";
defparam \in_wr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \Add0~4 (
	.dataa(\in_wr_ptr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[2] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[2]~q ),
	.prn(vcc));
defparam \in_wr_ptr[2] .is_wysiwyg = "true";
defparam \in_wr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add0~6 (
	.dataa(\in_wr_ptr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[3] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[3]~q ),
	.prn(vcc));
defparam \in_wr_ptr[3] .is_wysiwyg = "true";
defparam \in_wr_ptr[3] .power_up = "low";

cycloneive_lcell_comb \Add0~8 (
	.dataa(\in_wr_ptr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[4] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[4]~q ),
	.prn(vcc));
defparam \in_wr_ptr[4] .is_wysiwyg = "true";
defparam \in_wr_ptr[4] .power_up = "low";

cycloneive_lcell_comb \Add0~10 (
	.dataa(\in_wr_ptr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[5] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~10_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[5]~q ),
	.prn(vcc));
defparam \in_wr_ptr[5] .is_wysiwyg = "true";
defparam \in_wr_ptr[5] .power_up = "low";

cycloneive_lcell_comb \Add0~12 (
	.dataa(\in_wr_ptr[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[6] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[6]~q ),
	.prn(vcc));
defparam \in_wr_ptr[6] .is_wysiwyg = "true";
defparam \in_wr_ptr[6] .power_up = "low";

cycloneive_lcell_comb \Add0~14 (
	.dataa(\in_wr_ptr[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

dffeas \in_wr_ptr[7] (
	.clk(wire_pll7_clk_1),
	.d(\Add0~14_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_wr_ptr[7]~q ),
	.prn(vcc));
defparam \in_wr_ptr[7] .is_wysiwyg = "true";
defparam \in_wr_ptr[7] .power_up = "low";

cycloneive_lcell_comb \Add0~16 (
	.dataa(\in_wr_ptr[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout());
defparam \Add0~16 .lut_mask = 16'h5A5A;
defparam \Add0~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \next_in_rd_ptr[7]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\read_crosser|sync[8].u|dreg[1]~q ),
	.datad(\read_crosser|sync[7].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\next_in_rd_ptr[7]~0_combout ),
	.cout());
defparam \next_in_rd_ptr[7]~0 .lut_mask = 16'h0FF0;
defparam \next_in_rd_ptr[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_in_rd_ptr[3]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\next_in_rd_ptr[5]~2_combout ),
	.datad(\read_crosser|sync[4].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\next_in_rd_ptr[3]~3_combout ),
	.cout());
defparam \next_in_rd_ptr[3]~3 .lut_mask = 16'h0FF0;
defparam \next_in_rd_ptr[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_in_rd_ptr[0]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\next_in_rd_ptr[1]~5_combout ),
	.datad(\read_crosser|sync[1].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\next_in_rd_ptr[0]~6_combout ),
	.cout());
defparam \next_in_rd_ptr[0]~6 .lut_mask = 16'h0FF0;
defparam \next_in_rd_ptr[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_space_avail[0]~9 (
	.dataa(\Add0~0_combout ),
	.datab(\next_in_rd_ptr[0]~combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\in_space_avail[0]~9_combout ),
	.cout(\in_space_avail[0]~10 ));
defparam \in_space_avail[0]~9 .lut_mask = 16'h66DD;
defparam \in_space_avail[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_space_avail[1]~11 (
	.dataa(\Add0~2_combout ),
	.datab(\next_in_rd_ptr[0]~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[0]~10 ),
	.combout(\in_space_avail[1]~11_combout ),
	.cout(\in_space_avail[1]~12 ));
defparam \in_space_avail[1]~11 .lut_mask = 16'h96BF;
defparam \in_space_avail[1]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[2]~13 (
	.dataa(\Add0~4_combout ),
	.datab(\next_in_rd_ptr[1]~5_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[1]~12 ),
	.combout(\in_space_avail[2]~13_combout ),
	.cout(\in_space_avail[2]~14 ));
defparam \in_space_avail[2]~13 .lut_mask = 16'h96DF;
defparam \in_space_avail[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[3]~15 (
	.dataa(\Add0~6_combout ),
	.datab(\next_in_rd_ptr[3]~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[2]~14 ),
	.combout(\in_space_avail[3]~15_combout ),
	.cout(\in_space_avail[3]~16 ));
defparam \in_space_avail[3]~15 .lut_mask = 16'h96BF;
defparam \in_space_avail[3]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[4]~17 (
	.dataa(\Add0~8_combout ),
	.datab(\next_in_rd_ptr[3]~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[3]~16 ),
	.combout(\in_space_avail[4]~17_combout ),
	.cout(\in_space_avail[4]~18 ));
defparam \in_space_avail[4]~17 .lut_mask = 16'h96DF;
defparam \in_space_avail[4]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[5]~19 (
	.dataa(\Add0~10_combout ),
	.datab(\next_in_rd_ptr[5]~2_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[4]~18 ),
	.combout(\in_space_avail[5]~19_combout ),
	.cout(\in_space_avail[5]~20 ));
defparam \in_space_avail[5]~19 .lut_mask = 16'h96BF;
defparam \in_space_avail[5]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[6]~21 (
	.dataa(\Add0~12_combout ),
	.datab(\next_in_rd_ptr[5]~1_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[5]~20 ),
	.combout(\in_space_avail[6]~21_combout ),
	.cout(\in_space_avail[6]~22 ));
defparam \in_space_avail[6]~21 .lut_mask = 16'h96DF;
defparam \in_space_avail[6]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[7]~23 (
	.dataa(\Add0~14_combout ),
	.datab(\next_in_rd_ptr[7]~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\in_space_avail[6]~22 ),
	.combout(\in_space_avail[7]~23_combout ),
	.cout(\in_space_avail[7]~24 ));
defparam \in_space_avail[7]~23 .lut_mask = 16'h96BF;
defparam \in_space_avail[7]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \in_space_avail[8]~25 (
	.dataa(\Add0~16_combout ),
	.datab(\read_crosser|sync[8].u|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\in_space_avail[7]~24 ),
	.combout(\in_space_avail[8]~25_combout ),
	.cout());
defparam \in_space_avail[8]~25 .lut_mask = 16'h9696;
defparam \in_space_avail[8]~25 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[1] (
	.clk(clk_clk),
	.d(\Add1~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[1]~q ),
	.prn(vcc));
defparam \out_rd_ptr[1] .is_wysiwyg = "true";
defparam \out_rd_ptr[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\empty~q ),
	.datab(\out_rd_ptr[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
defparam \Add1~0 .lut_mask = 16'h66EE;
defparam \Add1~0 .sum_lutc_input = "datac";

dffeas \out_rd_ptr[0] (
	.clk(clk_clk),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[0]~q ),
	.prn(vcc));
defparam \out_rd_ptr[0] .is_wysiwyg = "true";
defparam \out_rd_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(\out_rd_ptr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Add1~0_combout ),
	.datad(\write_crosser|sync[0].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h0FF0;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\write_crosser|sync[5].u|dreg[1]~q ),
	.datab(\write_crosser|sync[6].u|dreg[1]~q ),
	.datac(\write_crosser|sync[7].u|dreg[1]~q ),
	.datad(\write_crosser|sync[8].u|dreg[1]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\write_crosser|sync[2].u|dreg[1]~q ),
	.datab(\write_crosser|sync[3].u|dreg[1]~q ),
	.datac(\write_crosser|sync[4].u|dreg[1]~q ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h6996;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\Add1~2_combout ),
	.datab(\Equal0~0_combout ),
	.datac(\write_crosser|sync[1].u|dreg[1]~q ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h6996;
defparam \Equal0~3 .sum_lutc_input = "datac";

dffeas \out_rd_ptr[8] (
	.clk(clk_clk),
	.d(\Add1~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[8]~q ),
	.prn(vcc));
defparam \out_rd_ptr[8] .is_wysiwyg = "true";
defparam \out_rd_ptr[8] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(\out_rd_ptr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
defparam \Add1~4 .lut_mask = 16'h5AAF;
defparam \Add1~4 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[2] (
	.clk(clk_clk),
	.d(\Add1~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[2]~q ),
	.prn(vcc));
defparam \out_rd_ptr[2] .is_wysiwyg = "true";
defparam \out_rd_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(\out_rd_ptr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[3] (
	.clk(clk_clk),
	.d(\Add1~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[3]~q ),
	.prn(vcc));
defparam \out_rd_ptr[3] .is_wysiwyg = "true";
defparam \out_rd_ptr[3] .power_up = "low";

cycloneive_lcell_comb \Add1~8 (
	.dataa(\out_rd_ptr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
defparam \Add1~8 .lut_mask = 16'h5AAF;
defparam \Add1~8 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[4] (
	.clk(clk_clk),
	.d(\Add1~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[4]~q ),
	.prn(vcc));
defparam \out_rd_ptr[4] .is_wysiwyg = "true";
defparam \out_rd_ptr[4] .power_up = "low";

cycloneive_lcell_comb \Add1~10 (
	.dataa(\out_rd_ptr[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
defparam \Add1~10 .lut_mask = 16'h5A5F;
defparam \Add1~10 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[5] (
	.clk(clk_clk),
	.d(\Add1~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[5]~q ),
	.prn(vcc));
defparam \out_rd_ptr[5] .is_wysiwyg = "true";
defparam \out_rd_ptr[5] .power_up = "low";

cycloneive_lcell_comb \Add1~12 (
	.dataa(\out_rd_ptr[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
defparam \Add1~12 .lut_mask = 16'h5AAF;
defparam \Add1~12 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[6] (
	.clk(clk_clk),
	.d(\Add1~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[6]~q ),
	.prn(vcc));
defparam \out_rd_ptr[6] .is_wysiwyg = "true";
defparam \out_rd_ptr[6] .power_up = "low";

cycloneive_lcell_comb \Add1~14 (
	.dataa(\out_rd_ptr[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
defparam \Add1~14 .lut_mask = 16'h5A5F;
defparam \Add1~14 .sum_lutc_input = "cin";

dffeas \out_rd_ptr[7] (
	.clk(clk_clk),
	.d(\Add1~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_rd_ptr[7]~q ),
	.prn(vcc));
defparam \out_rd_ptr[7] .is_wysiwyg = "true";
defparam \out_rd_ptr[7] .power_up = "low";

cycloneive_lcell_comb \Add1~16 (
	.dataa(\out_rd_ptr[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout());
defparam \Add1~16 .lut_mask = 16'h5A5A;
defparam \Add1~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\write_crosser|sync[8].u|dreg[1]~q ),
	.datab(\Add1~16_combout ),
	.datac(\write_crosser|sync[7].u|dreg[1]~q ),
	.datad(\Add1~14_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'h6996;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\Equal0~1_combout ),
	.datab(\Add1~10_combout ),
	.datac(\write_crosser|sync[4].u|dreg[1]~q ),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'h96FF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\write_crosser|sync[3].u|dreg[1]~q ),
	.datab(\Add1~6_combout ),
	.datac(\Add1~8_combout ),
	.datad(\Equal0~5_combout ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hB77B;
defparam \Equal0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~7 (
	.dataa(\write_crosser|sync[2].u|dreg[1]~q ),
	.datab(\Add1~4_combout ),
	.datac(\Add1~6_combout ),
	.datad(\Equal0~6_combout ),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'h6996;
defparam \Equal0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~8 (
	.dataa(\write_crosser|sync[6].u|dreg[1]~q ),
	.datab(\write_crosser|sync[7].u|dreg[1]~q ),
	.datac(\write_crosser|sync[8].u|dreg[1]~q ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'h6996;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~9 (
	.dataa(\Equal0~3_combout ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\Equal0~8_combout ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hFF7F;
defparam \Equal0~9 .sum_lutc_input = "datac";

dffeas empty(
	.clk(clk_clk),
	.d(\Equal0~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a0 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a0 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a1 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a1 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a2 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a2 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a3 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a3 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a4 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a4 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a5 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a5 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a6 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a6 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a7 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a7 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a8 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_8}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a8 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_first_bit_number = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_first_bit_number = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a9 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_9}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a9 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_first_bit_number = 9;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_first_bit_number = 9;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a10 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_10}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a10 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_first_bit_number = 10;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_first_bit_number = 10;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a11 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a11 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_first_bit_number = 11;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_first_bit_number = 11;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a12 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_12}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a12 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_first_bit_number = 12;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_first_bit_number = 12;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a13 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_13}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a13 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_first_bit_number = 13;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_first_bit_number = 13;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a14 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_14}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a14 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_first_bit_number = 14;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_first_bit_number = 14;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a15 (
	.portawe(\next_in_wr_ptr~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(wire_pll7_clk_1),
	.clk1(clk_clk),
	.ena0(\next_in_wr_ptr~0_combout ),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,av_readdata_pre_15}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\in_wr_ptr[7]~q ,\in_wr_ptr[6]~q ,\in_wr_ptr[5]~q ,\in_wr_ptr[4]~q ,\in_wr_ptr[3]~q ,\in_wr_ptr[2]~q ,\in_wr_ptr[1]~q ,\in_wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Add1~14_combout ,\Add1~12_combout ,\Add1~10_combout ,\Add1~8_combout ,\Add1~6_combout ,\Add1~4_combout ,\Add1~2_combout ,\Add1~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a15 .clk0_core_clock_enable = "ena0";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .logical_ram_name = "altera_avalon_mm_clock_crossing_bridge:clock_crossing_io|altera_avalon_dc_fifo:rsp_fifo|altsyncram:mem_rtl_0|altsyncram_e3d1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .mixed_port_feed_through_mode = "dont_care";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_first_bit_number = 15;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_first_bit_number = 15;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_last_address = 255;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_depth = 256;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_width = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_read_enable_clock = "clock1";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .ram_block_type = "auto";

endmodule

module usb_system_altera_dcfifo_synchronizer_bundle_2 (
	wire_pll7_clk_1,
	altera_reset_synchronizer_int_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	out_rd_ptr_gray_8,
	out_rd_ptr_gray_7,
	out_rd_ptr_gray_6,
	out_rd_ptr_gray_5,
	out_rd_ptr_gray_4,
	out_rd_ptr_gray_3,
	out_rd_ptr_gray_2,
	out_rd_ptr_gray_1,
	out_rd_ptr_gray_0)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
input 	altera_reset_synchronizer_int_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
input 	out_rd_ptr_gray_8;
input 	out_rd_ptr_gray_7;
input 	out_rd_ptr_gray_6;
input 	out_rd_ptr_gray_5;
input 	out_rd_ptr_gray_4;
input 	out_rd_ptr_gray_3;
input 	out_rd_ptr_gray_2;
input 	out_rd_ptr_gray_1;
input 	out_rd_ptr_gray_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_std_synchronizer_nocut_20 \sync[8].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_1),
	.din(out_rd_ptr_gray_8));

usb_system_altera_std_synchronizer_nocut_19 \sync[7].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_11),
	.din(out_rd_ptr_gray_7));

usb_system_altera_std_synchronizer_nocut_18 \sync[6].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_12),
	.din(out_rd_ptr_gray_6));

usb_system_altera_std_synchronizer_nocut_17 \sync[5].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_13),
	.din(out_rd_ptr_gray_5));

usb_system_altera_std_synchronizer_nocut_16 \sync[4].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_14),
	.din(out_rd_ptr_gray_4));

usb_system_altera_std_synchronizer_nocut_15 \sync[3].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_15),
	.din(out_rd_ptr_gray_3));

usb_system_altera_std_synchronizer_nocut_14 \sync[2].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_16),
	.din(out_rd_ptr_gray_2));

usb_system_altera_std_synchronizer_nocut_13 \sync[1].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_17),
	.din(out_rd_ptr_gray_1));

usb_system_altera_std_synchronizer_nocut_12 \sync[0].u (
	.clk(wire_pll7_clk_1),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_1(dreg_18),
	.din(out_rd_ptr_gray_0));

endmodule

module usb_system_altera_std_synchronizer_nocut_12 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_13 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_14 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_15 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_16 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_17 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_18 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_19 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_20 (
	clk,
	reset_n,
	dreg_1,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_1;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_dcfifo_synchronizer_bundle_3 (
	r_sync_rst,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	in_wr_ptr_gray_0,
	in_wr_ptr_gray_1,
	in_wr_ptr_gray_2,
	in_wr_ptr_gray_3,
	in_wr_ptr_gray_4,
	in_wr_ptr_gray_5,
	in_wr_ptr_gray_6,
	in_wr_ptr_gray_7,
	in_wr_ptr_gray_8,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
input 	in_wr_ptr_gray_0;
input 	in_wr_ptr_gray_1;
input 	in_wr_ptr_gray_2;
input 	in_wr_ptr_gray_3;
input 	in_wr_ptr_gray_4;
input 	in_wr_ptr_gray_5;
input 	in_wr_ptr_gray_6;
input 	in_wr_ptr_gray_7;
input 	in_wr_ptr_gray_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_std_synchronizer_nocut_29 \sync[8].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_18),
	.din(in_wr_ptr_gray_8),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_28 \sync[7].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_17),
	.din(in_wr_ptr_gray_7),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_27 \sync[6].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_16),
	.din(in_wr_ptr_gray_6),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_26 \sync[5].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_15),
	.din(in_wr_ptr_gray_5),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_25 \sync[4].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_14),
	.din(in_wr_ptr_gray_4),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_24 \sync[3].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_13),
	.din(in_wr_ptr_gray_3),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_23 \sync[2].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_12),
	.din(in_wr_ptr_gray_2),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_22 \sync[1].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_11),
	.din(in_wr_ptr_gray_1),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_nocut_21 \sync[0].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_1),
	.din(in_wr_ptr_gray_0),
	.clk(clk_clk));

endmodule

module usb_system_altera_std_synchronizer_nocut_21 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_22 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_23 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_24 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_25 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_26 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_27 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_28 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_nocut_29 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_irq_clock_crosser (
	r_sync_rst,
	dreg_1,
	oINT,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	dreg_1;
input 	oINT;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_std_synchronizer_bundle sync(
	.r_sync_rst(r_sync_rst),
	.dreg_1(dreg_1),
	.oINT(oINT),
	.clk_clk(clk_clk));

endmodule

module usb_system_altera_std_synchronizer_bundle (
	r_sync_rst,
	dreg_1,
	oINT,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	dreg_1;
input 	oINT;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_std_synchronizer \sync[0].u (
	.reset_n(r_sync_rst),
	.dreg_1(dreg_1),
	.din(oINT),
	.clk(clk_clk));

endmodule

module usb_system_altera_std_synchronizer (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module usb_system_altera_reset_controller (
	wire_pll7_clk_1,
	altera_reset_synchronizer_int_chain_out,
	resetrequest,
	merged_reset,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
output 	altera_reset_synchronizer_int_chain_out;
input 	resetrequest;
output 	merged_reset;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_reset_synchronizer_7 alt_rst_sync_uq1(
	.clk(wire_pll7_clk_1),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.merged_reset(merged_reset));

cycloneive_lcell_comb \merged_reset~0 (
	.dataa(resetrequest),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_reset_n),
	.cin(gnd),
	.combout(merged_reset),
	.cout());
defparam \merged_reset~0 .lut_mask = 16'hAAFF;
defparam \merged_reset~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_reset_controller_1 (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module usb_system_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module usb_system_altera_reset_controller_2 (
	r_sync_rst1,
	merged_reset,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
input 	merged_reset;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


usb_system_altera_reset_synchronizer_2 alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

usb_system_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.merged_reset(merged_reset),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 16'h5555;
defparam \altera_reset_synchronizer_int_chain[4]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.cout());
defparam \r_sync_rst_chain~1 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~1 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\altera_reset_synchronizer_int_chain[4]~q ),
	.datab(r_sync_rst1),
	.datac(gnd),
	.datad(\r_sync_rst_chain[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_reset_synchronizer_2 (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module usb_system_altera_reset_synchronizer_3 (
	merged_reset,
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	merged_reset;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module usb_system_altera_reset_controller_3 (
	wire_pll7_clk_0,
	altera_reset_synchronizer_int_chain_out,
	merged_reset)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_reset_synchronizer_5 alt_rst_sync_uq1(
	.clk(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.merged_reset(merged_reset));

endmodule

module usb_system_altera_reset_synchronizer_5 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	merged_reset)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module usb_system_altera_reset_synchronizer_7 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	merged_reset)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module usb_system_CY7C67200_IF (
	iCLK,
	HPI_ADDR_0,
	HPI_ADDR_1,
	HPI_RD_N1,
	HPI_WR_N1,
	HPI_CS_N1,
	iRST_N,
	out_payload_42,
	out_payload_43,
	av_read,
	av_write,
	TMP_DATA_0,
	TMP_DATA_1,
	TMP_DATA_2,
	TMP_DATA_3,
	TMP_DATA_4,
	TMP_DATA_5,
	TMP_DATA_6,
	TMP_DATA_7,
	TMP_DATA_8,
	TMP_DATA_9,
	TMP_DATA_10,
	TMP_DATA_11,
	TMP_DATA_12,
	TMP_DATA_13,
	TMP_DATA_14,
	TMP_DATA_15,
	iDATA,
	oDATA_0,
	oDATA_1,
	oDATA_2,
	oDATA_3,
	oDATA_4,
	oDATA_5,
	oDATA_6,
	oDATA_7,
	oDATA_8,
	oINT1,
	oDATA_9,
	oDATA_10,
	oDATA_11,
	oDATA_12,
	oDATA_13,
	oDATA_14,
	oDATA_15,
	av_begintransfer,
	usb_DATA_0,
	usb_DATA_1,
	usb_DATA_2,
	usb_DATA_3,
	usb_DATA_4,
	usb_DATA_5,
	usb_DATA_6,
	usb_DATA_7,
	usb_DATA_8,
	usb_DATA_9,
	usb_DATA_10,
	usb_DATA_11,
	usb_DATA_12,
	usb_DATA_13,
	usb_DATA_14,
	usb_DATA_15,
	usb_INT)/* synthesis synthesis_greybox=1 */;
input 	iCLK;
output 	HPI_ADDR_0;
output 	HPI_ADDR_1;
output 	HPI_RD_N1;
output 	HPI_WR_N1;
output 	HPI_CS_N1;
input 	iRST_N;
input 	out_payload_42;
input 	out_payload_43;
input 	av_read;
input 	av_write;
output 	TMP_DATA_0;
output 	TMP_DATA_1;
output 	TMP_DATA_2;
output 	TMP_DATA_3;
output 	TMP_DATA_4;
output 	TMP_DATA_5;
output 	TMP_DATA_6;
output 	TMP_DATA_7;
output 	TMP_DATA_8;
output 	TMP_DATA_9;
output 	TMP_DATA_10;
output 	TMP_DATA_11;
output 	TMP_DATA_12;
output 	TMP_DATA_13;
output 	TMP_DATA_14;
output 	TMP_DATA_15;
input 	[31:0] iDATA;
output 	oDATA_0;
output 	oDATA_1;
output 	oDATA_2;
output 	oDATA_3;
output 	oDATA_4;
output 	oDATA_5;
output 	oDATA_6;
output 	oDATA_7;
output 	oDATA_8;
output 	oINT1;
output 	oDATA_9;
output 	oDATA_10;
output 	oDATA_11;
output 	oDATA_12;
output 	oDATA_13;
output 	oDATA_14;
output 	oDATA_15;
input 	av_begintransfer;
input 	usb_DATA_0;
input 	usb_DATA_1;
input 	usb_DATA_2;
input 	usb_DATA_3;
input 	usb_DATA_4;
input 	usb_DATA_5;
input 	usb_DATA_6;
input 	usb_DATA_7;
input 	usb_DATA_8;
input 	usb_DATA_9;
input 	usb_DATA_10;
input 	usb_DATA_11;
input 	usb_DATA_12;
input 	usb_DATA_13;
input 	usb_DATA_14;
input 	usb_DATA_15;
input 	usb_INT;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \HPI_ADDR[0] (
	.clk(iCLK),
	.d(out_payload_42),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(HPI_ADDR_0),
	.prn(vcc));
defparam \HPI_ADDR[0] .is_wysiwyg = "true";
defparam \HPI_ADDR[0] .power_up = "low";

dffeas \HPI_ADDR[1] (
	.clk(iCLK),
	.d(out_payload_43),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(HPI_ADDR_1),
	.prn(vcc));
defparam \HPI_ADDR[1] .is_wysiwyg = "true";
defparam \HPI_ADDR[1] .power_up = "low";

dffeas HPI_RD_N(
	.clk(iCLK),
	.d(av_read),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(HPI_RD_N1),
	.prn(vcc));
defparam HPI_RD_N.is_wysiwyg = "true";
defparam HPI_RD_N.power_up = "low";

dffeas HPI_WR_N(
	.clk(iCLK),
	.d(av_write),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(HPI_WR_N1),
	.prn(vcc));
defparam HPI_WR_N.is_wysiwyg = "true";
defparam HPI_WR_N.power_up = "low";

dffeas HPI_CS_N(
	.clk(iCLK),
	.d(av_begintransfer),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(HPI_CS_N1),
	.prn(vcc));
defparam HPI_CS_N.is_wysiwyg = "true";
defparam HPI_CS_N.power_up = "low";

dffeas \TMP_DATA[0] (
	.clk(iCLK),
	.d(iDATA[0]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_0),
	.prn(vcc));
defparam \TMP_DATA[0] .is_wysiwyg = "true";
defparam \TMP_DATA[0] .power_up = "low";

dffeas \TMP_DATA[1] (
	.clk(iCLK),
	.d(iDATA[1]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_1),
	.prn(vcc));
defparam \TMP_DATA[1] .is_wysiwyg = "true";
defparam \TMP_DATA[1] .power_up = "low";

dffeas \TMP_DATA[2] (
	.clk(iCLK),
	.d(iDATA[2]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_2),
	.prn(vcc));
defparam \TMP_DATA[2] .is_wysiwyg = "true";
defparam \TMP_DATA[2] .power_up = "low";

dffeas \TMP_DATA[3] (
	.clk(iCLK),
	.d(iDATA[3]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_3),
	.prn(vcc));
defparam \TMP_DATA[3] .is_wysiwyg = "true";
defparam \TMP_DATA[3] .power_up = "low";

dffeas \TMP_DATA[4] (
	.clk(iCLK),
	.d(iDATA[4]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_4),
	.prn(vcc));
defparam \TMP_DATA[4] .is_wysiwyg = "true";
defparam \TMP_DATA[4] .power_up = "low";

dffeas \TMP_DATA[5] (
	.clk(iCLK),
	.d(iDATA[5]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_5),
	.prn(vcc));
defparam \TMP_DATA[5] .is_wysiwyg = "true";
defparam \TMP_DATA[5] .power_up = "low";

dffeas \TMP_DATA[6] (
	.clk(iCLK),
	.d(iDATA[6]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_6),
	.prn(vcc));
defparam \TMP_DATA[6] .is_wysiwyg = "true";
defparam \TMP_DATA[6] .power_up = "low";

dffeas \TMP_DATA[7] (
	.clk(iCLK),
	.d(iDATA[7]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_7),
	.prn(vcc));
defparam \TMP_DATA[7] .is_wysiwyg = "true";
defparam \TMP_DATA[7] .power_up = "low";

dffeas \TMP_DATA[8] (
	.clk(iCLK),
	.d(iDATA[8]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_8),
	.prn(vcc));
defparam \TMP_DATA[8] .is_wysiwyg = "true";
defparam \TMP_DATA[8] .power_up = "low";

dffeas \TMP_DATA[9] (
	.clk(iCLK),
	.d(iDATA[9]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_9),
	.prn(vcc));
defparam \TMP_DATA[9] .is_wysiwyg = "true";
defparam \TMP_DATA[9] .power_up = "low";

dffeas \TMP_DATA[10] (
	.clk(iCLK),
	.d(iDATA[10]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_10),
	.prn(vcc));
defparam \TMP_DATA[10] .is_wysiwyg = "true";
defparam \TMP_DATA[10] .power_up = "low";

dffeas \TMP_DATA[11] (
	.clk(iCLK),
	.d(iDATA[11]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_11),
	.prn(vcc));
defparam \TMP_DATA[11] .is_wysiwyg = "true";
defparam \TMP_DATA[11] .power_up = "low";

dffeas \TMP_DATA[12] (
	.clk(iCLK),
	.d(iDATA[12]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_12),
	.prn(vcc));
defparam \TMP_DATA[12] .is_wysiwyg = "true";
defparam \TMP_DATA[12] .power_up = "low";

dffeas \TMP_DATA[13] (
	.clk(iCLK),
	.d(iDATA[13]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_13),
	.prn(vcc));
defparam \TMP_DATA[13] .is_wysiwyg = "true";
defparam \TMP_DATA[13] .power_up = "low";

dffeas \TMP_DATA[14] (
	.clk(iCLK),
	.d(iDATA[14]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_14),
	.prn(vcc));
defparam \TMP_DATA[14] .is_wysiwyg = "true";
defparam \TMP_DATA[14] .power_up = "low";

dffeas \TMP_DATA[15] (
	.clk(iCLK),
	.d(iDATA[15]),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(TMP_DATA_15),
	.prn(vcc));
defparam \TMP_DATA[15] .is_wysiwyg = "true";
defparam \TMP_DATA[15] .power_up = "low";

dffeas \oDATA[0] (
	.clk(iCLK),
	.d(usb_DATA_0),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_0),
	.prn(vcc));
defparam \oDATA[0] .is_wysiwyg = "true";
defparam \oDATA[0] .power_up = "low";

dffeas \oDATA[1] (
	.clk(iCLK),
	.d(usb_DATA_1),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_1),
	.prn(vcc));
defparam \oDATA[1] .is_wysiwyg = "true";
defparam \oDATA[1] .power_up = "low";

dffeas \oDATA[2] (
	.clk(iCLK),
	.d(usb_DATA_2),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_2),
	.prn(vcc));
defparam \oDATA[2] .is_wysiwyg = "true";
defparam \oDATA[2] .power_up = "low";

dffeas \oDATA[3] (
	.clk(iCLK),
	.d(usb_DATA_3),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_3),
	.prn(vcc));
defparam \oDATA[3] .is_wysiwyg = "true";
defparam \oDATA[3] .power_up = "low";

dffeas \oDATA[4] (
	.clk(iCLK),
	.d(usb_DATA_4),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_4),
	.prn(vcc));
defparam \oDATA[4] .is_wysiwyg = "true";
defparam \oDATA[4] .power_up = "low";

dffeas \oDATA[5] (
	.clk(iCLK),
	.d(usb_DATA_5),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_5),
	.prn(vcc));
defparam \oDATA[5] .is_wysiwyg = "true";
defparam \oDATA[5] .power_up = "low";

dffeas \oDATA[6] (
	.clk(iCLK),
	.d(usb_DATA_6),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_6),
	.prn(vcc));
defparam \oDATA[6] .is_wysiwyg = "true";
defparam \oDATA[6] .power_up = "low";

dffeas \oDATA[7] (
	.clk(iCLK),
	.d(usb_DATA_7),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_7),
	.prn(vcc));
defparam \oDATA[7] .is_wysiwyg = "true";
defparam \oDATA[7] .power_up = "low";

dffeas \oDATA[8] (
	.clk(iCLK),
	.d(usb_DATA_8),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_8),
	.prn(vcc));
defparam \oDATA[8] .is_wysiwyg = "true";
defparam \oDATA[8] .power_up = "low";

dffeas oINT(
	.clk(iCLK),
	.d(usb_INT),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oINT1),
	.prn(vcc));
defparam oINT.is_wysiwyg = "true";
defparam oINT.power_up = "low";

dffeas \oDATA[9] (
	.clk(iCLK),
	.d(usb_DATA_9),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_9),
	.prn(vcc));
defparam \oDATA[9] .is_wysiwyg = "true";
defparam \oDATA[9] .power_up = "low";

dffeas \oDATA[10] (
	.clk(iCLK),
	.d(usb_DATA_10),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_10),
	.prn(vcc));
defparam \oDATA[10] .is_wysiwyg = "true";
defparam \oDATA[10] .power_up = "low";

dffeas \oDATA[11] (
	.clk(iCLK),
	.d(usb_DATA_11),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_11),
	.prn(vcc));
defparam \oDATA[11] .is_wysiwyg = "true";
defparam \oDATA[11] .power_up = "low";

dffeas \oDATA[12] (
	.clk(iCLK),
	.d(usb_DATA_12),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_12),
	.prn(vcc));
defparam \oDATA[12] .is_wysiwyg = "true";
defparam \oDATA[12] .power_up = "low";

dffeas \oDATA[13] (
	.clk(iCLK),
	.d(usb_DATA_13),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_13),
	.prn(vcc));
defparam \oDATA[13] .is_wysiwyg = "true";
defparam \oDATA[13] .power_up = "low";

dffeas \oDATA[14] (
	.clk(iCLK),
	.d(usb_DATA_14),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_14),
	.prn(vcc));
defparam \oDATA[14] .is_wysiwyg = "true";
defparam \oDATA[14] .power_up = "low";

dffeas \oDATA[15] (
	.clk(iCLK),
	.d(usb_DATA_15),
	.asdata(vcc),
	.clrn(iRST_N),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oDATA_15),
	.prn(vcc));
defparam \oDATA[15] .is_wysiwyg = "true";
defparam \oDATA[15] .power_up = "low";

endmodule

module usb_system_usb_system_all_switches (
	W_alu_result_2,
	W_alu_result_3,
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	clk_clk,
	all_switches_wire_export_0,
	all_switches_wire_export_1,
	all_switches_wire_export_2,
	all_switches_wire_export_3,
	all_switches_wire_export_4,
	all_switches_wire_export_5,
	all_switches_wire_export_6,
	all_switches_wire_export_7,
	all_switches_wire_export_8,
	all_switches_wire_export_9,
	all_switches_wire_export_10,
	all_switches_wire_export_11,
	all_switches_wire_export_12,
	all_switches_wire_export_13,
	all_switches_wire_export_14,
	all_switches_wire_export_15,
	all_switches_wire_export_16,
	all_switches_wire_export_17)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
input 	clk_clk;
input 	all_switches_wire_export_0;
input 	all_switches_wire_export_1;
input 	all_switches_wire_export_2;
input 	all_switches_wire_export_3;
input 	all_switches_wire_export_4;
input 	all_switches_wire_export_5;
input 	all_switches_wire_export_6;
input 	all_switches_wire_export_7;
input 	all_switches_wire_export_8;
input 	all_switches_wire_export_9;
input 	all_switches_wire_export_10;
input 	all_switches_wire_export_11;
input 	all_switches_wire_export_12;
input 	all_switches_wire_export_13;
input 	all_switches_wire_export_14;
input 	all_switches_wire_export_15;
input 	all_switches_wire_export_16;
input 	all_switches_wire_export_17;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;
wire \read_mux_out[8]~combout ;
wire \read_mux_out[9]~combout ;
wire \read_mux_out[10]~combout ;
wire \read_mux_out[11]~combout ;
wire \read_mux_out[12]~combout ;
wire \read_mux_out[13]~combout ;
wire \read_mux_out[14]~combout ;
wire \read_mux_out[15]~combout ;
wire \read_mux_out[16]~combout ;
wire \read_mux_out[17]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\read_mux_out[8]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\read_mux_out[9]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\read_mux_out[10]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\read_mux_out[11]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\read_mux_out[12]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\read_mux_out[13]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\read_mux_out[14]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\read_mux_out[15]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\read_mux_out[16]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\read_mux_out[17]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

cycloneive_lcell_comb \read_mux_out[0] (
	.dataa(all_switches_wire_export_0),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[0]~combout ),
	.cout());
defparam \read_mux_out[0] .lut_mask = 16'hAFFF;
defparam \read_mux_out[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[1] (
	.dataa(all_switches_wire_export_1),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[1]~combout ),
	.cout());
defparam \read_mux_out[1] .lut_mask = 16'hAFFF;
defparam \read_mux_out[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[2] (
	.dataa(all_switches_wire_export_2),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[2]~combout ),
	.cout());
defparam \read_mux_out[2] .lut_mask = 16'hAFFF;
defparam \read_mux_out[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[3] (
	.dataa(all_switches_wire_export_3),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[3]~combout ),
	.cout());
defparam \read_mux_out[3] .lut_mask = 16'hAFFF;
defparam \read_mux_out[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[4] (
	.dataa(all_switches_wire_export_4),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[4]~combout ),
	.cout());
defparam \read_mux_out[4] .lut_mask = 16'hAFFF;
defparam \read_mux_out[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[5] (
	.dataa(all_switches_wire_export_5),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[5]~combout ),
	.cout());
defparam \read_mux_out[5] .lut_mask = 16'hAFFF;
defparam \read_mux_out[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[6] (
	.dataa(all_switches_wire_export_6),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[6]~combout ),
	.cout());
defparam \read_mux_out[6] .lut_mask = 16'hAFFF;
defparam \read_mux_out[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[7] (
	.dataa(all_switches_wire_export_7),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[7]~combout ),
	.cout());
defparam \read_mux_out[7] .lut_mask = 16'hAFFF;
defparam \read_mux_out[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[8] (
	.dataa(all_switches_wire_export_8),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[8]~combout ),
	.cout());
defparam \read_mux_out[8] .lut_mask = 16'hAFFF;
defparam \read_mux_out[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[9] (
	.dataa(all_switches_wire_export_9),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[9]~combout ),
	.cout());
defparam \read_mux_out[9] .lut_mask = 16'hAFFF;
defparam \read_mux_out[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[10] (
	.dataa(all_switches_wire_export_10),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[10]~combout ),
	.cout());
defparam \read_mux_out[10] .lut_mask = 16'hAFFF;
defparam \read_mux_out[10] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[11] (
	.dataa(all_switches_wire_export_11),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[11]~combout ),
	.cout());
defparam \read_mux_out[11] .lut_mask = 16'hAFFF;
defparam \read_mux_out[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[12] (
	.dataa(all_switches_wire_export_12),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[12]~combout ),
	.cout());
defparam \read_mux_out[12] .lut_mask = 16'hAFFF;
defparam \read_mux_out[12] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[13] (
	.dataa(all_switches_wire_export_13),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[13]~combout ),
	.cout());
defparam \read_mux_out[13] .lut_mask = 16'hAFFF;
defparam \read_mux_out[13] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[14] (
	.dataa(all_switches_wire_export_14),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[14]~combout ),
	.cout());
defparam \read_mux_out[14] .lut_mask = 16'hAFFF;
defparam \read_mux_out[14] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[15] (
	.dataa(all_switches_wire_export_15),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[15]~combout ),
	.cout());
defparam \read_mux_out[15] .lut_mask = 16'hAFFF;
defparam \read_mux_out[15] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[16] (
	.dataa(all_switches_wire_export_16),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[16]~combout ),
	.cout());
defparam \read_mux_out[16] .lut_mask = 16'hAFFF;
defparam \read_mux_out[16] .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_mux_out[17] (
	.dataa(all_switches_wire_export_17),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\read_mux_out[17]~combout ),
	.cout());
defparam \read_mux_out[17] .lut_mask = 16'hAFFF;
defparam \read_mux_out[17] .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_clocks (
	wire_pll7_clk_0,
	wire_pll7_clk_1,
	d_writedata_0,
	reset,
	d_writedata_1,
	mem_used_1,
	WideOr1,
	src_data_38,
	mem,
	src_data_39,
	mem1,
	readdata_0,
	readdata_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	wire_pll7_clk_0;
output 	wire_pll7_clk_1;
input 	d_writedata_0;
input 	reset;
input 	d_writedata_1;
input 	mem_used_1;
input 	WideOr1;
input 	src_data_38;
input 	mem;
input 	src_data_39;
input 	mem1;
output 	readdata_0;
output 	readdata_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \stdsync2|dffpipe3|dffe6a[0]~q ;
wire \sd1|locked~combout ;
wire \readdata[0]~0_combout ;
wire \w_reset~0_combout ;
wire \w_reset~1_combout ;
wire \prev_reset~q ;
wire \pfdena_reg~0_combout ;
wire \pfdena_reg~q ;


usb_system_usb_system_clocks_altpll_pqa2 sd1(
	.clk({clk_unconnected_wire_4,clk_unconnected_wire_3,clk_unconnected_wire_2,wire_pll7_clk_1,wire_pll7_clk_0}),
	.areset(\prev_reset~q ),
	.locked1(\sd1|locked~combout ),
	.inclk({gnd,clk_clk}));

usb_system_usb_system_clocks_stdsync_sv6 stdsync2(
	.r_sync_rst(reset),
	.dffe6a_0(\stdsync2|dffpipe3|dffe6a[0]~q ),
	.locked(\sd1|locked~combout ),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \readdata[0]~1 (
	.dataa(\readdata[0]~0_combout ),
	.datab(\prev_reset~q ),
	.datac(\stdsync2|dffpipe3|dffe6a[0]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0]~1 .lut_mask = 16'hFAFC;
defparam \readdata[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1]~2 (
	.dataa(\readdata[0]~0_combout ),
	.datab(gnd),
	.datac(src_data_38),
	.datad(\pfdena_reg~q ),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1]~2 .lut_mask = 16'hAFFF;
defparam \readdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~0 (
	.dataa(WideOr1),
	.datab(mem1),
	.datac(mem_used_1),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\readdata[0]~0_combout ),
	.cout());
defparam \readdata[0]~0 .lut_mask = 16'hEFFF;
defparam \readdata[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \w_reset~0 (
	.dataa(WideOr1),
	.datab(src_data_38),
	.datac(mem),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\w_reset~0_combout ),
	.cout());
defparam \w_reset~0 .lut_mask = 16'hFEFF;
defparam \w_reset~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \w_reset~1 (
	.dataa(d_writedata_0),
	.datab(\w_reset~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\w_reset~1_combout ),
	.cout());
defparam \w_reset~1 .lut_mask = 16'hEEEE;
defparam \w_reset~1 .sum_lutc_input = "datac";

dffeas prev_reset(
	.clk(clk_clk),
	.d(\w_reset~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prev_reset~q ),
	.prn(vcc));
defparam prev_reset.is_wysiwyg = "true";
defparam prev_reset.power_up = "low";

cycloneive_lcell_comb \pfdena_reg~0 (
	.dataa(d_writedata_1),
	.datab(\w_reset~0_combout ),
	.datac(gnd),
	.datad(\pfdena_reg~q ),
	.cin(gnd),
	.combout(\pfdena_reg~0_combout ),
	.cout());
defparam \pfdena_reg~0 .lut_mask = 16'hDD11;
defparam \pfdena_reg~0 .sum_lutc_input = "datac";

dffeas pfdena_reg(
	.clk(clk_clk),
	.d(\pfdena_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pfdena_reg~q ),
	.prn(vcc));
defparam pfdena_reg.is_wysiwyg = "true";
defparam pfdena_reg.power_up = "low";

endmodule

module usb_system_usb_system_clocks_altpll_pqa2 (
	clk,
	areset,
	locked1,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	[4:0] clk;
input 	areset;
output 	locked1;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wire_pll7_clk[2] ;
wire \wire_pll7_clk[3] ;
wire \wire_pll7_clk[4] ;
wire wire_pll7_locked;
wire wire_pll7_fbout;
wire \pll_lock_sync~q ;

wire [4:0] pll7_CLK_bus;

assign clk[0] = pll7_CLK_bus[0];
assign clk[1] = pll7_CLK_bus[1];
assign \wire_pll7_clk[2]  = pll7_CLK_bus[2];
assign \wire_pll7_clk[3]  = pll7_CLK_bus[3];
assign \wire_pll7_clk[4]  = pll7_CLK_bus[4];

cycloneive_pll pll7(
	.areset(areset),
	.pfdena(vcc),
	.fbin(wire_pll7_fbout),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scandata(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect(3'b000),
	.phasedone(),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(wire_pll7_locked),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(wire_pll7_fbout),
	.clk(pll7_CLK_bus),
	.clkbad());
defparam pll7.auto_settings = "false";
defparam pll7.bandwidth_type = "auto";
defparam pll7.c0_high = 10;
defparam pll7.c0_initial = 1;
defparam pll7.c0_low = 10;
defparam pll7.c0_mode = "even";
defparam pll7.c0_ph = 0;
defparam pll7.c1_high = 50;
defparam pll7.c1_initial = 4;
defparam pll7.c1_low = 50;
defparam pll7.c1_mode = "even";
defparam pll7.c1_ph = 0;
defparam pll7.c1_use_casc_in = "off";
defparam pll7.c2_high = 1;
defparam pll7.c2_initial = 1;
defparam pll7.c2_low = 1;
defparam pll7.c2_mode = "bypass";
defparam pll7.c2_ph = 0;
defparam pll7.c2_use_casc_in = "off";
defparam pll7.c3_high = 1;
defparam pll7.c3_initial = 1;
defparam pll7.c3_low = 1;
defparam pll7.c3_mode = "bypass";
defparam pll7.c3_ph = 0;
defparam pll7.c3_use_casc_in = "off";
defparam pll7.c4_high = 1;
defparam pll7.c4_initial = 1;
defparam pll7.c4_low = 1;
defparam pll7.c4_mode = "bypass";
defparam pll7.c4_ph = 0;
defparam pll7.c4_use_casc_in = "off";
defparam pll7.charge_pump_current_bits = 2;
defparam pll7.clk0_counter = "c0";
defparam pll7.clk0_divide_by = 1;
defparam pll7.clk0_duty_cycle = 50;
defparam pll7.clk0_multiply_by = 1;
defparam pll7.clk0_phase_shift = "-3000";
defparam pll7.clk1_counter = "c1";
defparam pll7.clk1_divide_by = 5;
defparam pll7.clk1_duty_cycle = 50;
defparam pll7.clk1_multiply_by = 1;
defparam pll7.clk1_phase_shift = "0";
defparam pll7.clk2_counter = "unused";
defparam pll7.clk2_divide_by = 0;
defparam pll7.clk2_duty_cycle = 50;
defparam pll7.clk2_multiply_by = 0;
defparam pll7.clk2_phase_shift = "0";
defparam pll7.clk3_counter = "unused";
defparam pll7.clk3_divide_by = 0;
defparam pll7.clk3_duty_cycle = 50;
defparam pll7.clk3_multiply_by = 0;
defparam pll7.clk3_phase_shift = "0";
defparam pll7.clk4_counter = "unused";
defparam pll7.clk4_divide_by = 0;
defparam pll7.clk4_duty_cycle = 50;
defparam pll7.clk4_multiply_by = 0;
defparam pll7.clk4_phase_shift = "0";
defparam pll7.compensate_clock = "clock0";
defparam pll7.inclk0_input_frequency = 20000;
defparam pll7.inclk1_input_frequency = 0;
defparam pll7.loop_filter_c_bits = 2;
defparam pll7.loop_filter_r_bits = 1;
defparam pll7.m = 20;
defparam pll7.m_initial = 4;
defparam pll7.m_ph = 0;
defparam pll7.n = 1;
defparam pll7.operation_mode = "normal";
defparam pll7.pfd_max = 0;
defparam pll7.pfd_min = 0;
defparam pll7.self_reset_on_loss_lock = "off";
defparam pll7.simulation_type = "timing";
defparam pll7.switch_over_type = "auto";
defparam pll7.vco_center = 0;
defparam pll7.vco_divide_by = 0;
defparam pll7.vco_frequency_control = "auto";
defparam pll7.vco_max = 0;
defparam pll7.vco_min = 0;
defparam pll7.vco_multiply_by = 0;
defparam pll7.vco_phase_shift_step = 0;
defparam pll7.vco_post_scale = 1;

cycloneive_lcell_comb locked(
	.dataa(wire_pll7_locked),
	.datab(\pll_lock_sync~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(locked1),
	.cout());
defparam locked.lut_mask = 16'hEEEE;
defparam locked.sum_lutc_input = "datac";

dffeas pll_lock_sync(
	.clk(wire_pll7_locked),
	.d(vcc),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_lock_sync~q ),
	.prn(vcc));
defparam pll_lock_sync.is_wysiwyg = "true";
defparam pll_lock_sync.power_up = "low";

endmodule

module usb_system_usb_system_clocks_stdsync_sv6 (
	r_sync_rst,
	dffe6a_0,
	locked,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	dffe6a_0;
input 	locked;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_usb_system_clocks_dffpipe_l2c dffpipe3(
	.clrn(r_sync_rst),
	.dffe6a_0(dffe6a_0),
	.d({locked}),
	.clock(clk_clk));

endmodule

module usb_system_usb_system_clocks_dffpipe_l2c (
	clrn,
	dffe6a_0,
	d,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clrn;
output 	dffe6a_0;
input 	[0:0] d;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe4a[0]~q ;
wire \dffe5a[0]~q ;


dffeas \dffe6a[0] (
	.clk(clock),
	.d(\dffe5a[0]~q ),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe6a_0),
	.prn(vcc));
defparam \dffe6a[0] .is_wysiwyg = "true";
defparam \dffe6a[0] .power_up = "low";

dffeas \dffe4a[0] (
	.clk(clock),
	.d(d[0]),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe4a[0]~q ),
	.prn(vcc));
defparam \dffe4a[0] .is_wysiwyg = "true";
defparam \dffe4a[0] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock),
	.d(\dffe4a[0]~q ),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe5a[0]~q ),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

endmodule

module usb_system_usb_system_cpu (
	sr_0,
	W_alu_result_7,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_8,
	W_alu_result_6,
	W_alu_result_24,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_5,
	readdata_6,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	debug_reset_request,
	d_read,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	out_valid,
	src0_valid,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	mem_86_0,
	mem_68_0,
	src0_valid1,
	read_latency_shift_reg_04,
	read_latency_shift_reg_05,
	WideOr1,
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	src0_valid2,
	mem_67_04,
	mem_67_05,
	mem_67_06,
	mem_67_07,
	mem_67_08,
	out_valid1,
	out_data_buffer_67,
	av_ld_getting_data,
	debug_mem_slave_waitrequest,
	mem_used_1,
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_5,
	F_pc_6,
	F_pc_4,
	F_pc_1,
	F_pc_3,
	i_read,
	F_pc_2,
	av_waitrequest,
	F_pc_0,
	WideOr11,
	local_read,
	src1_valid,
	src_payload,
	out_valid2,
	src_payload1,
	WideOr12,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	hbreak_enabled,
	out_data_buffer_0,
	av_readdata_pre_0,
	av_readdata_pre_01,
	out_data_buffer_1,
	av_readdata_pre_1,
	av_readdata_pre_11,
	out_data_buffer_2,
	av_readdata_pre_2,
	av_readdata_pre_30,
	src_payload2,
	av_readdata_pre_3,
	out_data_buffer_4,
	av_readdata_pre_4,
	src_data_0,
	out_data_buffer_22,
	av_readdata_pre_22,
	av_readdata_pre_23,
	out_data_buffer_23,
	out_data_buffer_24,
	av_readdata_pre_24,
	av_readdata_pre_25,
	out_data_buffer_25,
	out_data_buffer_26,
	av_readdata_pre_26,
	out_data_buffer_11,
	av_readdata_pre_111,
	out_data_buffer_13,
	av_readdata_pre_13,
	src_payload3,
	av_readdata_pre_16,
	av_readdata_pre_12,
	out_data_buffer_12,
	out_data_buffer_5,
	av_readdata_pre_5,
	out_data_buffer_14,
	av_readdata_pre_14,
	out_data_buffer_15,
	av_readdata_pre_15,
	av_readdata_pre_10,
	out_data_buffer_10,
	out_data_buffer_9,
	av_readdata_pre_9,
	out_data_buffer_8,
	av_readdata_pre_8,
	out_data_buffer_7,
	av_readdata_pre_7,
	out_data_buffer_6,
	av_readdata_pre_6,
	src_payload4,
	av_readdata_pre_20,
	out_data_buffer_18,
	av_readdata_pre_18,
	out_data_buffer_19,
	av_readdata_pre_19,
	out_data_buffer_17,
	av_readdata_pre_17,
	src_payload5,
	av_readdata_pre_21,
	av_readdata_pre_27,
	out_data_buffer_27,
	out_data_buffer_28,
	av_readdata_pre_28,
	av_readdata_pre_31,
	out_data_buffer_31,
	out_data_buffer_30,
	av_readdata_pre_301,
	av_readdata_pre_29,
	out_data_buffer_29,
	mem,
	src_data_46,
	src_data_1,
	src_payload6,
	src_data_2,
	src_data_3,
	src_data_31,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	src_data_8,
	dreg_1,
	av_readdata_9,
	av_readdata_8,
	readdata_4,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	r_early_rst,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_14,
	readdata_15,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_20,
	readdata_18,
	readdata_19,
	readdata_17,
	src_payload7,
	readdata_21,
	src_payload8,
	readdata_27,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	out_data_buffer_241,
	readdata_28,
	out_data_buffer_281,
	out_data_buffer_271,
	readdata_31,
	out_data_buffer_261,
	readdata_30,
	out_data_buffer_251,
	readdata_29,
	src_payload13,
	src_payload14,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	out_data_buffer_311,
	out_data_buffer_301,
	out_data_buffer_291,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_34,
	src_payload22,
	src_payload23,
	src_payload24,
	src_data_35,
	src_payload25,
	src_payload26,
	src_payload27,
	src_data_33,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_data_21,
	src_data_47,
	src_data_51,
	src_data_61,
	src_data_71,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_7;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_23;
output 	W_alu_result_22;
output 	W_alu_result_8;
output 	W_alu_result_6;
output 	W_alu_result_24;
output 	W_alu_result_21;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_28;
output 	W_alu_result_27;
output 	W_alu_result_26;
output 	W_alu_result_25;
output 	W_alu_result_4;
output 	W_alu_result_5;
output 	W_alu_result_2;
output 	W_alu_result_3;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_5;
output 	readdata_6;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_10;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
output 	debug_reset_request;
output 	d_read;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	out_valid;
input 	src0_valid;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	mem_86_0;
input 	mem_68_0;
input 	src0_valid1;
input 	read_latency_shift_reg_04;
input 	read_latency_shift_reg_05;
input 	WideOr1;
input 	mem_67_0;
input 	mem_67_01;
input 	mem_67_02;
input 	mem_67_03;
input 	src0_valid2;
input 	mem_67_04;
input 	mem_67_05;
input 	mem_67_06;
input 	mem_67_07;
input 	mem_67_08;
input 	out_valid1;
input 	out_data_buffer_67;
output 	av_ld_getting_data;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
output 	F_pc_26;
output 	F_pc_25;
output 	F_pc_24;
output 	F_pc_23;
output 	F_pc_22;
output 	F_pc_21;
output 	F_pc_20;
output 	F_pc_19;
output 	F_pc_18;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_9;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_5;
output 	F_pc_6;
output 	F_pc_4;
output 	F_pc_1;
output 	F_pc_3;
output 	i_read;
output 	F_pc_2;
input 	av_waitrequest;
output 	F_pc_0;
input 	WideOr11;
input 	local_read;
input 	src1_valid;
input 	src_payload;
input 	out_valid2;
input 	src_payload1;
input 	WideOr12;
input 	av_readdatavalid;
input 	av_readdatavalid1;
input 	av_readdatavalid2;
output 	hbreak_enabled;
input 	out_data_buffer_0;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	out_data_buffer_1;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	out_data_buffer_2;
input 	av_readdata_pre_2;
input 	av_readdata_pre_30;
input 	src_payload2;
input 	av_readdata_pre_3;
input 	out_data_buffer_4;
input 	av_readdata_pre_4;
input 	src_data_0;
input 	out_data_buffer_22;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	out_data_buffer_23;
input 	out_data_buffer_24;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	out_data_buffer_25;
input 	out_data_buffer_26;
input 	av_readdata_pre_26;
input 	out_data_buffer_11;
input 	av_readdata_pre_111;
input 	out_data_buffer_13;
input 	av_readdata_pre_13;
input 	src_payload3;
input 	av_readdata_pre_16;
input 	av_readdata_pre_12;
input 	out_data_buffer_12;
input 	out_data_buffer_5;
input 	av_readdata_pre_5;
input 	out_data_buffer_14;
input 	av_readdata_pre_14;
input 	out_data_buffer_15;
input 	av_readdata_pre_15;
input 	av_readdata_pre_10;
input 	out_data_buffer_10;
input 	out_data_buffer_9;
input 	av_readdata_pre_9;
input 	out_data_buffer_8;
input 	av_readdata_pre_8;
input 	out_data_buffer_7;
input 	av_readdata_pre_7;
input 	out_data_buffer_6;
input 	av_readdata_pre_6;
input 	src_payload4;
input 	av_readdata_pre_20;
input 	out_data_buffer_18;
input 	av_readdata_pre_18;
input 	out_data_buffer_19;
input 	av_readdata_pre_19;
input 	out_data_buffer_17;
input 	av_readdata_pre_17;
input 	src_payload5;
input 	av_readdata_pre_21;
input 	av_readdata_pre_27;
input 	out_data_buffer_27;
input 	out_data_buffer_28;
input 	av_readdata_pre_28;
input 	av_readdata_pre_31;
input 	out_data_buffer_31;
input 	out_data_buffer_30;
input 	av_readdata_pre_301;
input 	av_readdata_pre_29;
input 	out_data_buffer_29;
input 	mem;
input 	src_data_46;
input 	src_data_1;
input 	src_payload6;
input 	src_data_2;
input 	src_data_3;
input 	src_data_31;
input 	src_data_4;
input 	src_data_5;
input 	src_data_6;
input 	src_data_7;
input 	src_data_8;
input 	dreg_1;
input 	av_readdata_9;
input 	av_readdata_8;
output 	readdata_4;
input 	src_data_9;
input 	src_data_10;
input 	src_data_11;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_data_17;
output 	d_byteenable_0;
output 	d_byteenable_1;
output 	d_byteenable_2;
output 	d_byteenable_3;
input 	r_early_rst;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_20;
output 	readdata_18;
output 	readdata_19;
output 	readdata_17;
input 	src_payload7;
output 	readdata_21;
input 	src_payload8;
output 	readdata_27;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	out_data_buffer_241;
output 	readdata_28;
input 	out_data_buffer_281;
input 	out_data_buffer_271;
output 	readdata_31;
input 	out_data_buffer_261;
output 	readdata_30;
input 	out_data_buffer_251;
output 	readdata_29;
input 	src_payload13;
input 	src_payload14;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
input 	out_data_buffer_311;
input 	out_data_buffer_301;
input 	out_data_buffer_291;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
output 	d_writedata_18;
output 	d_writedata_19;
output 	d_writedata_20;
output 	d_writedata_21;
output 	d_writedata_22;
output 	d_writedata_23;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_data_34;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_data_35;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_data_33;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	src_payload44;
input 	src_payload45;
input 	src_data_21;
input 	src_data_47;
input 	src_data_51;
input 	src_data_61;
input 	src_data_71;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_usb_system_cpu_cpu cpu(
	.sr_0(sr_0),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.readdata_5(readdata_5),
	.readdata_6(readdata_6),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_write1(d_write),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.debug_reset_request(debug_reset_request),
	.d_read1(d_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.out_valid(out_valid),
	.src0_valid(src0_valid),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.read_latency_shift_reg_03(read_latency_shift_reg_03),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_04(read_latency_shift_reg_04),
	.read_latency_shift_reg_05(read_latency_shift_reg_05),
	.WideOr1(WideOr1),
	.mem_67_0(mem_67_0),
	.mem_67_01(mem_67_01),
	.mem_67_02(mem_67_02),
	.mem_67_03(mem_67_03),
	.src0_valid2(src0_valid2),
	.mem_67_04(mem_67_04),
	.mem_67_05(mem_67_05),
	.mem_67_06(mem_67_06),
	.mem_67_07(mem_67_07),
	.mem_67_08(mem_67_08),
	.out_valid1(out_valid1),
	.out_data_buffer_67(out_data_buffer_67),
	.av_ld_getting_data(av_ld_getting_data),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.F_pc_26(F_pc_26),
	.F_pc_25(F_pc_25),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_4(F_pc_4),
	.F_pc_1(F_pc_1),
	.F_pc_3(F_pc_3),
	.i_read1(i_read),
	.F_pc_2(F_pc_2),
	.av_waitrequest(av_waitrequest),
	.F_pc_0(F_pc_0),
	.WideOr11(WideOr11),
	.local_read(local_read),
	.src1_valid(src1_valid),
	.src_payload(src_payload),
	.out_valid2(out_valid2),
	.src_payload1(src_payload1),
	.WideOr12(WideOr12),
	.av_readdatavalid(av_readdatavalid),
	.av_readdatavalid1(av_readdatavalid1),
	.av_readdatavalid2(av_readdatavalid2),
	.hbreak_enabled1(hbreak_enabled),
	.out_data_buffer_0(out_data_buffer_0),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_01(av_readdata_pre_01),
	.out_data_buffer_1(out_data_buffer_1),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_11(av_readdata_pre_11),
	.out_data_buffer_2(out_data_buffer_2),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_30(av_readdata_pre_30),
	.src_payload2(src_payload2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.out_data_buffer_4(out_data_buffer_4),
	.av_readdata_pre_4(av_readdata_pre_4),
	.src_data_0(src_data_0),
	.out_data_buffer_22(out_data_buffer_22),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_24(out_data_buffer_24),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_26(out_data_buffer_26),
	.av_readdata_pre_26(av_readdata_pre_26),
	.out_data_buffer_11(out_data_buffer_11),
	.av_readdata_pre_111(av_readdata_pre_111),
	.out_data_buffer_13(out_data_buffer_13),
	.av_readdata_pre_13(av_readdata_pre_13),
	.src_payload3(src_payload3),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.av_readdata_pre_5(av_readdata_pre_5),
	.out_data_buffer_14(out_data_buffer_14),
	.av_readdata_pre_14(av_readdata_pre_14),
	.out_data_buffer_15(out_data_buffer_15),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_10(av_readdata_pre_10),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.av_readdata_pre_9(av_readdata_pre_9),
	.out_data_buffer_8(out_data_buffer_8),
	.av_readdata_pre_8(av_readdata_pre_8),
	.out_data_buffer_7(out_data_buffer_7),
	.av_readdata_pre_7(av_readdata_pre_7),
	.out_data_buffer_6(out_data_buffer_6),
	.av_readdata_pre_6(av_readdata_pre_6),
	.src_payload4(src_payload4),
	.av_readdata_pre_20(av_readdata_pre_20),
	.out_data_buffer_18(out_data_buffer_18),
	.av_readdata_pre_18(av_readdata_pre_18),
	.out_data_buffer_19(out_data_buffer_19),
	.av_readdata_pre_19(av_readdata_pre_19),
	.out_data_buffer_17(out_data_buffer_17),
	.av_readdata_pre_17(av_readdata_pre_17),
	.src_payload5(src_payload5),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_27(av_readdata_pre_27),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_28(out_data_buffer_28),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_31(av_readdata_pre_31),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.av_readdata_pre_301(av_readdata_pre_301),
	.av_readdata_pre_29(av_readdata_pre_29),
	.out_data_buffer_29(out_data_buffer_29),
	.mem(mem),
	.src_data_46(src_data_46),
	.src_data_1(src_data_1),
	.src_payload6(src_payload6),
	.src_data_2(src_data_2),
	.src_data_3(src_data_3),
	.src_data_31(src_data_31),
	.src_data_4(src_data_4),
	.src_data_5(src_data_5),
	.src_data_6(src_data_6),
	.src_data_7(src_data_7),
	.src_data_8(src_data_8),
	.dreg_1(dreg_1),
	.av_readdata_9(av_readdata_9),
	.av_readdata_8(av_readdata_8),
	.readdata_4(readdata_4),
	.src_data_9(src_data_9),
	.src_data_10(src_data_10),
	.src_data_11(src_data_11),
	.src_data_12(src_data_12),
	.src_data_13(src_data_13),
	.src_data_14(src_data_14),
	.src_data_15(src_data_15),
	.src_data_16(src_data_16),
	.src_data_17(src_data_17),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.r_early_rst(r_early_rst),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_11(readdata_11),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_20(readdata_20),
	.readdata_18(readdata_18),
	.readdata_19(readdata_19),
	.readdata_17(readdata_17),
	.src_payload7(src_payload7),
	.readdata_21(readdata_21),
	.src_payload8(src_payload8),
	.readdata_27(readdata_27),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.out_data_buffer_241(out_data_buffer_241),
	.readdata_28(readdata_28),
	.out_data_buffer_281(out_data_buffer_281),
	.out_data_buffer_271(out_data_buffer_271),
	.readdata_31(readdata_31),
	.out_data_buffer_261(out_data_buffer_261),
	.readdata_30(readdata_30),
	.out_data_buffer_251(out_data_buffer_251),
	.readdata_29(readdata_29),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.out_data_buffer_311(out_data_buffer_311),
	.out_data_buffer_301(out_data_buffer_301),
	.out_data_buffer_291(out_data_buffer_291),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_data_34(src_data_34),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_data_35(src_data_35),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_data_33(src_data_33),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.src_payload33(src_payload33),
	.src_payload34(src_payload34),
	.src_payload35(src_payload35),
	.src_payload36(src_payload36),
	.src_payload37(src_payload37),
	.src_payload38(src_payload38),
	.src_payload39(src_payload39),
	.src_payload40(src_payload40),
	.src_payload41(src_payload41),
	.src_payload42(src_payload42),
	.src_payload43(src_payload43),
	.src_payload44(src_payload44),
	.src_payload45(src_payload45),
	.src_data_21(src_data_21),
	.src_data_47(src_data_47),
	.src_data_51(src_data_51),
	.src_data_61(src_data_61),
	.src_data_71(src_data_71),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module usb_system_usb_system_cpu_cpu (
	sr_0,
	W_alu_result_7,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_8,
	W_alu_result_6,
	W_alu_result_24,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_5,
	readdata_6,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	debug_reset_request,
	d_read1,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	out_valid,
	src0_valid,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	mem_86_0,
	mem_68_0,
	src0_valid1,
	read_latency_shift_reg_04,
	read_latency_shift_reg_05,
	WideOr1,
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	src0_valid2,
	mem_67_04,
	mem_67_05,
	mem_67_06,
	mem_67_07,
	mem_67_08,
	out_valid1,
	out_data_buffer_67,
	av_ld_getting_data,
	debug_mem_slave_waitrequest,
	mem_used_1,
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_5,
	F_pc_6,
	F_pc_4,
	F_pc_1,
	F_pc_3,
	i_read1,
	F_pc_2,
	av_waitrequest,
	F_pc_0,
	WideOr11,
	local_read,
	src1_valid,
	src_payload,
	out_valid2,
	src_payload1,
	WideOr12,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	hbreak_enabled1,
	out_data_buffer_0,
	av_readdata_pre_0,
	av_readdata_pre_01,
	out_data_buffer_1,
	av_readdata_pre_1,
	av_readdata_pre_11,
	out_data_buffer_2,
	av_readdata_pre_2,
	av_readdata_pre_30,
	src_payload2,
	av_readdata_pre_3,
	out_data_buffer_4,
	av_readdata_pre_4,
	src_data_0,
	out_data_buffer_22,
	av_readdata_pre_22,
	av_readdata_pre_23,
	out_data_buffer_23,
	out_data_buffer_24,
	av_readdata_pre_24,
	av_readdata_pre_25,
	out_data_buffer_25,
	out_data_buffer_26,
	av_readdata_pre_26,
	out_data_buffer_11,
	av_readdata_pre_111,
	out_data_buffer_13,
	av_readdata_pre_13,
	src_payload3,
	av_readdata_pre_16,
	av_readdata_pre_12,
	out_data_buffer_12,
	out_data_buffer_5,
	av_readdata_pre_5,
	out_data_buffer_14,
	av_readdata_pre_14,
	out_data_buffer_15,
	av_readdata_pre_15,
	av_readdata_pre_10,
	out_data_buffer_10,
	out_data_buffer_9,
	av_readdata_pre_9,
	out_data_buffer_8,
	av_readdata_pre_8,
	out_data_buffer_7,
	av_readdata_pre_7,
	out_data_buffer_6,
	av_readdata_pre_6,
	src_payload4,
	av_readdata_pre_20,
	out_data_buffer_18,
	av_readdata_pre_18,
	out_data_buffer_19,
	av_readdata_pre_19,
	out_data_buffer_17,
	av_readdata_pre_17,
	src_payload5,
	av_readdata_pre_21,
	av_readdata_pre_27,
	out_data_buffer_27,
	out_data_buffer_28,
	av_readdata_pre_28,
	av_readdata_pre_31,
	out_data_buffer_31,
	out_data_buffer_30,
	av_readdata_pre_301,
	av_readdata_pre_29,
	out_data_buffer_29,
	mem,
	src_data_46,
	src_data_1,
	src_payload6,
	src_data_2,
	src_data_3,
	src_data_31,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	src_data_8,
	dreg_1,
	av_readdata_9,
	av_readdata_8,
	readdata_4,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	r_early_rst,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_14,
	readdata_15,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_20,
	readdata_18,
	readdata_19,
	readdata_17,
	src_payload7,
	readdata_21,
	src_payload8,
	readdata_27,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	out_data_buffer_241,
	readdata_28,
	out_data_buffer_281,
	out_data_buffer_271,
	readdata_31,
	out_data_buffer_261,
	readdata_30,
	out_data_buffer_251,
	readdata_29,
	src_payload13,
	src_payload14,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	out_data_buffer_311,
	out_data_buffer_301,
	out_data_buffer_291,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_34,
	src_payload22,
	src_payload23,
	src_payload24,
	src_data_35,
	src_payload25,
	src_payload26,
	src_payload27,
	src_data_33,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_data_21,
	src_data_47,
	src_data_51,
	src_data_61,
	src_data_71,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_7;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_12;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_23;
output 	W_alu_result_22;
output 	W_alu_result_8;
output 	W_alu_result_6;
output 	W_alu_result_24;
output 	W_alu_result_21;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_28;
output 	W_alu_result_27;
output 	W_alu_result_26;
output 	W_alu_result_25;
output 	W_alu_result_4;
output 	W_alu_result_5;
output 	W_alu_result_2;
output 	W_alu_result_3;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_5;
output 	readdata_6;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write1;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_10;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
output 	debug_reset_request;
output 	d_read1;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	out_valid;
input 	src0_valid;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	mem_86_0;
input 	mem_68_0;
input 	src0_valid1;
input 	read_latency_shift_reg_04;
input 	read_latency_shift_reg_05;
input 	WideOr1;
input 	mem_67_0;
input 	mem_67_01;
input 	mem_67_02;
input 	mem_67_03;
input 	src0_valid2;
input 	mem_67_04;
input 	mem_67_05;
input 	mem_67_06;
input 	mem_67_07;
input 	mem_67_08;
input 	out_valid1;
input 	out_data_buffer_67;
output 	av_ld_getting_data;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
output 	F_pc_26;
output 	F_pc_25;
output 	F_pc_24;
output 	F_pc_23;
output 	F_pc_22;
output 	F_pc_21;
output 	F_pc_20;
output 	F_pc_19;
output 	F_pc_18;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_9;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_5;
output 	F_pc_6;
output 	F_pc_4;
output 	F_pc_1;
output 	F_pc_3;
output 	i_read1;
output 	F_pc_2;
input 	av_waitrequest;
output 	F_pc_0;
input 	WideOr11;
input 	local_read;
input 	src1_valid;
input 	src_payload;
input 	out_valid2;
input 	src_payload1;
input 	WideOr12;
input 	av_readdatavalid;
input 	av_readdatavalid1;
input 	av_readdatavalid2;
output 	hbreak_enabled1;
input 	out_data_buffer_0;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	out_data_buffer_1;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	out_data_buffer_2;
input 	av_readdata_pre_2;
input 	av_readdata_pre_30;
input 	src_payload2;
input 	av_readdata_pre_3;
input 	out_data_buffer_4;
input 	av_readdata_pre_4;
input 	src_data_0;
input 	out_data_buffer_22;
input 	av_readdata_pre_22;
input 	av_readdata_pre_23;
input 	out_data_buffer_23;
input 	out_data_buffer_24;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	out_data_buffer_25;
input 	out_data_buffer_26;
input 	av_readdata_pre_26;
input 	out_data_buffer_11;
input 	av_readdata_pre_111;
input 	out_data_buffer_13;
input 	av_readdata_pre_13;
input 	src_payload3;
input 	av_readdata_pre_16;
input 	av_readdata_pre_12;
input 	out_data_buffer_12;
input 	out_data_buffer_5;
input 	av_readdata_pre_5;
input 	out_data_buffer_14;
input 	av_readdata_pre_14;
input 	out_data_buffer_15;
input 	av_readdata_pre_15;
input 	av_readdata_pre_10;
input 	out_data_buffer_10;
input 	out_data_buffer_9;
input 	av_readdata_pre_9;
input 	out_data_buffer_8;
input 	av_readdata_pre_8;
input 	out_data_buffer_7;
input 	av_readdata_pre_7;
input 	out_data_buffer_6;
input 	av_readdata_pre_6;
input 	src_payload4;
input 	av_readdata_pre_20;
input 	out_data_buffer_18;
input 	av_readdata_pre_18;
input 	out_data_buffer_19;
input 	av_readdata_pre_19;
input 	out_data_buffer_17;
input 	av_readdata_pre_17;
input 	src_payload5;
input 	av_readdata_pre_21;
input 	av_readdata_pre_27;
input 	out_data_buffer_27;
input 	out_data_buffer_28;
input 	av_readdata_pre_28;
input 	av_readdata_pre_31;
input 	out_data_buffer_31;
input 	out_data_buffer_30;
input 	av_readdata_pre_301;
input 	av_readdata_pre_29;
input 	out_data_buffer_29;
input 	mem;
input 	src_data_46;
input 	src_data_1;
input 	src_payload6;
input 	src_data_2;
input 	src_data_3;
input 	src_data_31;
input 	src_data_4;
input 	src_data_5;
input 	src_data_6;
input 	src_data_7;
input 	src_data_8;
input 	dreg_1;
input 	av_readdata_9;
input 	av_readdata_8;
output 	readdata_4;
input 	src_data_9;
input 	src_data_10;
input 	src_data_11;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_data_17;
output 	d_byteenable_0;
output 	d_byteenable_1;
output 	d_byteenable_2;
output 	d_byteenable_3;
input 	r_early_rst;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_20;
output 	readdata_18;
output 	readdata_19;
output 	readdata_17;
input 	src_payload7;
output 	readdata_21;
input 	src_payload8;
output 	readdata_27;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	out_data_buffer_241;
output 	readdata_28;
input 	out_data_buffer_281;
input 	out_data_buffer_271;
output 	readdata_31;
input 	out_data_buffer_261;
output 	readdata_30;
input 	out_data_buffer_251;
output 	readdata_29;
input 	src_payload13;
input 	src_payload14;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
input 	out_data_buffer_311;
input 	out_data_buffer_301;
input 	out_data_buffer_291;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
output 	d_writedata_18;
output 	d_writedata_19;
output 	d_writedata_20;
output 	d_writedata_21;
output 	d_writedata_22;
output 	d_writedata_23;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_data_34;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_data_35;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_data_33;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	src_payload44;
input 	src_payload45;
input 	src_data_21;
input 	src_data_47;
input 	src_data_51;
input 	src_data_61;
input 	src_data_71;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \W_alu_result[0]~q ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \W_alu_result[1]~q ;
wire \av_ld_byte1_data[0]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_oci_debug|jtag_break~q ;
wire \av_ld_byte1_data[1]~q ;
wire \av_ld_byte1_data[2]~q ;
wire \av_ld_byte1_data[3]~q ;
wire \av_ld_byte1_data[4]~q ;
wire \av_ld_byte1_data[5]~q ;
wire \av_ld_byte1_data[6]~q ;
wire \av_ld_byte1_data[7]~q ;
wire \av_ld_byte2_data[0]~q ;
wire \av_ld_byte2_data[1]~q ;
wire \Add1~92_combout ;
wire \Add1~94_combout ;
wire \Add1~96_combout ;
wire \W_alu_result[0]~27_combout ;
wire \av_ld_byte2_data[2]~q ;
wire \av_ld_byte2_data[7]~q ;
wire \av_ld_byte2_data[6]~q ;
wire \av_ld_byte2_data[5]~q ;
wire \av_ld_byte2_data[4]~q ;
wire \av_ld_byte2_data[3]~q ;
wire \W_alu_result[1]~28_combout ;
wire \av_ld_byte1_data[0]~0_combout ;
wire \av_ld_byte1_data[1]~1_combout ;
wire \av_ld_byte1_data[2]~2_combout ;
wire \av_ld_byte1_data[3]~3_combout ;
wire \av_ld_byte1_data[4]~4_combout ;
wire \av_ld_byte1_data[5]~5_combout ;
wire \av_ld_byte1_data[6]~6_combout ;
wire \av_ld_byte1_data[7]~7_combout ;
wire \av_ld_byte2_data[0]~0_combout ;
wire \av_ld_byte2_data[1]~1_combout ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \av_ld_byte2_data[2]~4_combout ;
wire \av_ld_byte2_data[7]~2_combout ;
wire \av_ld_byte2_data[6]~3_combout ;
wire \av_ld_byte2_data[5]~7_combout ;
wire \av_ld_byte2_data[4]~6_combout ;
wire \av_ld_byte2_data[3]~5_combout ;
wire \W_alu_result[31]~q ;
wire \W_alu_result[29]~q ;
wire \W_alu_result[30]~q ;
wire \W_alu_result[31]~29_combout ;
wire \W_alu_result[29]~30_combout ;
wire \W_alu_result[30]~31_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \av_ld_byte0_data[0]~q ;
wire \W_rf_wr_data[0]~0_combout ;
wire \W_control_rd_data[0]~q ;
wire \W_rf_wr_data[0]~1_combout ;
wire \W_rf_wr_data[0]~2_combout ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \av_ld_byte0_data[1]~q ;
wire \W_rf_wr_data[1]~3_combout ;
wire \av_ld_byte0_data[2]~q ;
wire \W_rf_wr_data[2]~4_combout ;
wire \av_ld_byte0_data[3]~q ;
wire \W_rf_wr_data[3]~5_combout ;
wire \av_ld_byte0_data[4]~q ;
wire \W_rf_wr_data[4]~6_combout ;
wire \av_ld_byte0_data[5]~q ;
wire \W_control_rd_data[5]~q ;
wire \W_rf_wr_data[5]~7_combout ;
wire \W_rf_wr_data[5]~8_combout ;
wire \av_ld_byte0_data[6]~q ;
wire \W_control_rd_data[6]~q ;
wire \W_rf_wr_data[6]~9_combout ;
wire \W_rf_wr_data[6]~10_combout ;
wire \av_ld_byte0_data[7]~q ;
wire \W_rf_wr_data[7]~11_combout ;
wire \W_rf_wr_data[8]~12_combout ;
wire \W_rf_wr_data[9]~13_combout ;
wire \W_rf_wr_data[10]~14_combout ;
wire \W_rf_wr_data[11]~15_combout ;
wire \W_rf_wr_data[12]~16_combout ;
wire \W_rf_wr_data[13]~17_combout ;
wire \W_rf_wr_data[14]~18_combout ;
wire \W_rf_wr_data[15]~19_combout ;
wire \W_rf_wr_data[16]~20_combout ;
wire \W_rf_wr_data[17]~21_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~1_combout ;
wire \Equal0~14_combout ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_dst_regnum[0]~1_combout ;
wire \D_dst_regnum[0]~2_combout ;
wire \D_dst_regnum[0]~3_combout ;
wire \D_dst_regnum[0]~12_combout ;
wire \D_dst_regnum[0]~13_combout ;
wire \D_dst_regnum[2]~14_combout ;
wire \D_dst_regnum[3]~15_combout ;
wire \D_dst_regnum[4]~16_combout ;
wire \Equal0~18_combout ;
wire \D_dst_regnum[1]~17_combout ;
wire \D_dst_regnum[1]~18_combout ;
wire \D_wr_dst_reg~2_combout ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_rshift8~1_combout ;
wire \av_ld_byte0_data[4]~0_combout ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_control_rd_data[0]~1_combout ;
wire \D_ctrl_ld_signed~1_combout ;
wire \W_rf_wr_data[18]~22_combout ;
wire \W_rf_wr_data[23]~23_combout ;
wire \W_rf_wr_data[22]~24_combout ;
wire \W_rf_wr_data[21]~25_combout ;
wire \W_rf_wr_data[20]~26_combout ;
wire \W_rf_wr_data[19]~27_combout ;
wire \av_ld_byte3_data[0]~q ;
wire \W_rf_wr_data[24]~28_combout ;
wire \av_ld_byte3_data[4]~q ;
wire \W_rf_wr_data[28]~29_combout ;
wire \av_ld_byte3_data[3]~q ;
wire \W_rf_wr_data[27]~30_combout ;
wire \av_ld_byte3_data[2]~q ;
wire \W_rf_wr_data[26]~31_combout ;
wire \av_ld_byte3_data[1]~q ;
wire \W_rf_wr_data[25]~32_combout ;
wire \av_ld_byte0_data_nxt[2]~4_combout ;
wire \av_ld_byte0_data_nxt[3]~5_combout ;
wire \av_ld_byte0_data_nxt[4]~6_combout ;
wire \av_ld_byte0_data_nxt[5]~7_combout ;
wire \E_control_rd_data[5]~2_combout ;
wire \E_control_rd_data[5]~3_combout ;
wire \av_ld_byte0_data_nxt[6]~8_combout ;
wire \E_control_rd_data[6]~4_combout ;
wire \av_ld_byte0_data_nxt[7]~9_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[6]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[5]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \av_ld_byte3_data[7]~q ;
wire \av_ld_byte3_data[6]~q ;
wire \av_ld_byte3_data[5]~q ;
wire \av_ld_byte3_data_nxt~0_combout ;
wire \av_ld_byte3_data_nxt~1_combout ;
wire \av_ld_byte3_data_nxt~2_combout ;
wire \av_ld_byte3_data_nxt~3_combout ;
wire \av_ld_byte3_data_nxt~4_combout ;
wire \av_ld_byte3_data_nxt~5_combout ;
wire \av_ld_byte3_data_nxt~6_combout ;
wire \av_ld_byte3_data_nxt~7_combout ;
wire \av_ld_byte3_data_nxt~8_combout ;
wire \av_ld_byte3_data_nxt~9_combout ;
wire \W_rf_wr_data[31]~33_combout ;
wire \W_rf_wr_data[29]~34_combout ;
wire \W_rf_wr_data[30]~35_combout ;
wire \av_ld_byte3_data_nxt~10_combout ;
wire \av_ld_byte3_data_nxt~11_combout ;
wire \av_ld_byte3_data_nxt~12_combout ;
wire \av_ld_byte3_data_nxt~13_combout ;
wire \av_ld_byte3_data_nxt~14_combout ;
wire \av_ld_byte3_data_nxt~15_combout ;
wire \av_ld_byte0_data_nxt[0]~10_combout ;
wire \av_ld_byte0_data_nxt[1]~11_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \F_iw[11]~25_combout ;
wire \F_iw[10]~37_combout ;
wire \F_iw[10]~38_combout ;
wire \D_iw[10]~q ;
wire \F_iw[4]~13_combout ;
wire \F_iw[4]~14_combout ;
wire \D_iw[4]~q ;
wire \F_iw[1]~8_combout ;
wire \F_iw[1]~9_combout ;
wire \D_iw[1]~q ;
wire \F_iw[0]~6_combout ;
wire \F_iw[0]~7_combout ;
wire \D_iw[0]~q ;
wire \F_iw[3]~12_combout ;
wire \D_iw[3]~q ;
wire \F_iw[2]~10_combout ;
wire \F_iw[2]~11_combout ;
wire \D_iw[2]~q ;
wire \Equal0~2_combout ;
wire \F_iw[5]~32_combout ;
wire \F_iw[5]~33_combout ;
wire \D_iw[5]~q ;
wire \Equal0~7_combout ;
wire \F_iw[15]~35_combout ;
wire \F_iw[15]~36_combout ;
wire \D_iw[15]~q ;
wire \E_new_inst~q ;
wire \D_ctrl_st~0_combout ;
wire \R_ctrl_st~q ;
wire \W_valid~3_combout ;
wire \W_valid~2_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \F_iw[14]~34_combout ;
wire \F_iw[14]~64_combout ;
wire \D_iw[14]~q ;
wire \D_op_opx_rsv63~0_combout ;
wire \F_iw[13]~27_combout ;
wire \F_iw[13]~28_combout ;
wire \D_iw[13]~q ;
wire \F_iw[16]~29_combout ;
wire \D_iw[16]~q ;
wire \F_iw[12]~30_combout ;
wire \F_iw[12]~31_combout ;
wire \D_iw[12]~q ;
wire \Equal62~4_combout ;
wire \Equal62~5_combout ;
wire \Equal62~6_combout ;
wire \D_ctrl_shift_rot~0_combout ;
wire \Equal62~7_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_shift_rot~3_combout ;
wire \R_ctrl_shift_rot~q ;
wire \E_shift_rot_cnt[0]~5_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~1_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \Equal0~12_combout ;
wire \D_ctrl_alu_force_xor~14_combout ;
wire \Equal0~17_combout ;
wire \Equal0~11_combout ;
wire \D_ctrl_exception~2_combout ;
wire \Equal62~14_combout ;
wire \Equal62~9_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal62~13_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \Equal0~16_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \D_ctrl_force_src2_zero~3_combout ;
wire \Equal0~3_combout ;
wire \D_op_opx_rsv00~0_combout ;
wire \Equal62~2_combout ;
wire \D_dst_regnum[0]~20_combout ;
wire \Equal62~10_combout ;
wire \Equal62~11_combout ;
wire \D_op_opx_rsv17~0_combout ;
wire \D_dst_regnum[0]~5_combout ;
wire \Equal62~8_combout ;
wire \D_op_cmpge~0_combout ;
wire \D_dst_regnum[0]~4_combout ;
wire \D_dst_regnum[0]~21_combout ;
wire \Equal0~15_combout ;
wire \D_dst_regnum[0]~6_combout ;
wire \Equal62~12_combout ;
wire \D_dst_regnum[0]~7_combout ;
wire \Equal62~1_combout ;
wire \Equal62~3_combout ;
wire \D_dst_regnum[0]~8_combout ;
wire \D_dst_regnum[0]~9_combout ;
wire \D_dst_regnum[0]~10_combout ;
wire \D_dst_regnum[0]~11_combout ;
wire \Equal0~4_combout ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_force_src2_zero~4_combout ;
wire \Equal0~19_combout ;
wire \D_ctrl_force_src2_zero~5_combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_force_src2_zero~6_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \R_src2_lo[2]~3_combout ;
wire \F_iw[6]~45_combout ;
wire \F_iw[6]~46_combout ;
wire \D_iw[6]~q ;
wire \D_dst_regnum[0]~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~5_combout ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~1_combout ;
wire \D_ctrl_b_is_dst~2_combout ;
wire \Equal0~13_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \R_ctrl_br_nxt~1_combout ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \E_src2[3]~16_combout ;
wire \R_src2_lo[0]~8_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~q ;
wire \E_shift_rot_cnt[0]~6 ;
wire \E_shift_rot_cnt[1]~7_combout ;
wire \F_iw[7]~43_combout ;
wire \F_iw[7]~44_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~7_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \E_shift_rot_cnt[1]~8 ;
wire \E_shift_rot_cnt[2]~9_combout ;
wire \F_iw[8]~41_combout ;
wire \F_iw[8]~42_combout ;
wire \D_iw[8]~q ;
wire \R_src2_lo[2]~6_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \E_stall~0_combout ;
wire \E_shift_rot_cnt[2]~10 ;
wire \E_shift_rot_cnt[3]~11_combout ;
wire \F_iw[9]~39_combout ;
wire \F_iw[9]~40_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~5_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_shift_rot_cnt[3]~12 ;
wire \E_shift_rot_cnt[4]~13_combout ;
wire \R_src2_lo[4]~4_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~1_combout ;
wire \E_stall~2_combout ;
wire \D_ctrl_ld_signed~0_combout ;
wire \D_ctrl_ld~2_combout ;
wire \D_ctrl_ld~3_combout ;
wire \R_ctrl_ld~q ;
wire \av_ld_getting_data~0_combout ;
wire \av_ld_getting_data~1_combout ;
wire \av_ld_getting_data~2_combout ;
wire \av_ld_getting_data~3_combout ;
wire \av_ld_getting_data~4_combout ;
wire \av_ld_getting_data~5_combout ;
wire \av_ld_getting_data~7_combout ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \av_ld_aligning_data~q ;
wire \av_ld_align_cycle_nxt[0]~0_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \D_ctrl_mem16~0_combout ;
wire \D_ctrl_mem16~1_combout ;
wire \av_ld_align_cycle_nxt[1]~1_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \E_stall~3_combout ;
wire \E_stall~4_combout ;
wire \E_valid_from_R~3_combout ;
wire \E_valid_from_R~2_combout ;
wire \E_valid_from_R~q ;
wire \D_ctrl_jmp_direct~1_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_src1~10_combout ;
wire \E_src1[6]~24_combout ;
wire \F_pc_plus_one[0]~1 ;
wire \F_pc_plus_one[1]~3 ;
wire \F_pc_plus_one[2]~5 ;
wire \F_pc_plus_one[3]~7 ;
wire \F_pc_plus_one[4]~8_combout ;
wire \R_ctrl_br~q ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_retaddr~4_combout ;
wire \D_ctrl_retaddr~5_combout ;
wire \Equal0~9_combout ;
wire \D_ctrl_retaddr~6_combout ;
wire \D_ctrl_retaddr~7_combout ;
wire \D_ctrl_retaddr~8_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~11_combout ;
wire \E_src1[6]~q ;
wire \D_op_wrctl~combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \W_ienable_reg_nxt~0_combout ;
wire \W_ienable_reg_nxt~1_combout ;
wire \W_ienable_reg[6]~q ;
wire \W_ipending_reg_nxt[6]~0_combout ;
wire \W_ipending_reg[6]~q ;
wire \E_src1[5]~25_combout ;
wire \F_pc_plus_one[3]~6_combout ;
wire \E_src1[5]~q ;
wire \W_ienable_reg[5]~q ;
wire \W_ipending_reg_nxt[5]~1_combout ;
wire \W_ipending_reg[5]~q ;
wire \R_src1[0]~13_combout ;
wire \E_src1[0]~q ;
wire \E_wrctl_estatus~0_combout ;
wire \D_ctrl_exception~4_combout ;
wire \D_dst_regnum[0]~19_combout ;
wire \D_ctrl_exception~5_combout ;
wire \D_ctrl_exception~6_combout ;
wire \D_ctrl_exception~0_combout ;
wire \D_ctrl_exception~1_combout ;
wire \D_ctrl_exception~3_combout ;
wire \D_ctrl_exception~7_combout ;
wire \R_ctrl_exception~q ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \W_estatus_reg_inst_nxt~1_combout ;
wire \W_estatus_reg~q ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \D_ctrl_break~0_combout ;
wire \R_ctrl_break~q ;
wire \W_bstatus_reg_inst_nxt~1_combout ;
wire \W_bstatus_reg~q ;
wire \E_wrctl_status~0_combout ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \D_op_eret~combout ;
wire \F_pc_sel_nxt.10~1_combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_status_reg_pie~q ;
wire \D_iw[5]~0_combout ;
wire \D_iw[5]~1_combout ;
wire \F_iw[11]~26_combout ;
wire \D_iw[11]~q ;
wire \Equal62~0_combout ;
wire \Equal0~5_combout ;
wire \D_ctrl_alu_subtract~8_combout ;
wire \D_ctrl_alu_subtract~9_combout ;
wire \D_ctrl_alu_subtract~5_combout ;
wire \D_ctrl_alu_subtract~10_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \E_src2[12]~15_combout ;
wire \R_src2_lo[7]~0_combout ;
wire \E_src2[7]~q ;
wire \Add1~0_combout ;
wire \E_src1[7]~23_combout ;
wire \F_pc_plus_one[4]~9 ;
wire \F_pc_plus_one[5]~10_combout ;
wire \E_src1[7]~q ;
wire \R_src2_lo[6]~1_combout ;
wire \E_src2[6]~q ;
wire \Add1~1_combout ;
wire \R_src2_lo[5]~2_combout ;
wire \E_src2[5]~q ;
wire \Add1~2_combout ;
wire \Add1~3_combout ;
wire \E_src1[4]~26_combout ;
wire \F_pc_plus_one[2]~4_combout ;
wire \E_src1[4]~q ;
wire \Add1~4_combout ;
wire \E_src1[3]~8_combout ;
wire \F_pc_plus_one[1]~2_combout ;
wire \E_src1[3]~q ;
wire \Add1~5_combout ;
wire \E_src1[2]~7_combout ;
wire \F_pc_plus_one[0]~0_combout ;
wire \E_src1[2]~q ;
wire \Add1~6_combout ;
wire \R_src1[1]~12_combout ;
wire \E_src1[1]~q ;
wire \Add1~7_combout ;
wire \Add1~9_cout ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~24_combout ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~10_combout ;
wire \D_ctrl_alu_force_xor~11_combout ;
wire \D_ctrl_alu_force_xor~13_combout ;
wire \D_ctrl_alu_force_xor~12_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[7]~0_combout ;
wire \Equal0~8_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~combout ;
wire \R_ctrl_logic~q ;
wire \W_alu_result[7]~23_combout ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \E_shift_rot_result_nxt[6]~14_combout ;
wire \E_shift_rot_result[6]~q ;
wire \E_shift_rot_result_nxt[5]~24_combout ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[4]~23_combout ;
wire \E_shift_rot_result[4]~q ;
wire \E_shift_rot_result_nxt[3]~26_combout ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[2]~25_combout ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[1]~28_combout ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[0]~29_combout ;
wire \E_shift_rot_result[0]~q ;
wire \R_ctrl_rot_right_nxt~0_combout ;
wire \R_ctrl_rot_right~q ;
wire \D_ctrl_shift_logical~1_combout ;
wire \D_ctrl_shift_logical~2_combout ;
wire \R_ctrl_shift_logical~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[31]~31_combout ;
wire \R_src1[31]~14_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_result_nxt[30]~30_combout ;
wire \R_src1[30]~16_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[29]~27_combout ;
wire \R_src1[29]~15_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[28]~19_combout ;
wire \E_src1[28]~0_combout ;
wire \F_pc_plus_one[5]~11 ;
wire \F_pc_plus_one[6]~13 ;
wire \F_pc_plus_one[7]~15 ;
wire \F_pc_plus_one[8]~17 ;
wire \F_pc_plus_one[9]~19 ;
wire \F_pc_plus_one[10]~21 ;
wire \F_pc_plus_one[11]~23 ;
wire \F_pc_plus_one[12]~25 ;
wire \F_pc_plus_one[13]~27 ;
wire \F_pc_plus_one[14]~29 ;
wire \F_pc_plus_one[15]~31 ;
wire \F_pc_plus_one[16]~33 ;
wire \F_pc_plus_one[17]~35 ;
wire \F_pc_plus_one[18]~37 ;
wire \F_pc_plus_one[19]~39 ;
wire \F_pc_plus_one[20]~41 ;
wire \F_pc_plus_one[21]~43 ;
wire \F_pc_plus_one[22]~45 ;
wire \F_pc_plus_one[23]~47 ;
wire \F_pc_plus_one[24]~49 ;
wire \F_pc_plus_one[25]~51 ;
wire \F_pc_plus_one[26]~52_combout ;
wire \E_src1[28]~q ;
wire \E_shift_rot_result[28]~q ;
wire \E_shift_rot_result_nxt[27]~20_combout ;
wire \F_iw[31]~58_combout ;
wire \F_iw[31]~59_combout ;
wire \D_iw[31]~q ;
wire \E_src1[27]~1_combout ;
wire \F_pc_plus_one[25]~50_combout ;
wire \E_src1[27]~q ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[26]~21_combout ;
wire \F_iw[30]~60_combout ;
wire \F_iw[30]~61_combout ;
wire \D_iw[30]~q ;
wire \E_src1[26]~2_combout ;
wire \F_pc_plus_one[24]~48_combout ;
wire \E_src1[26]~q ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[25]~22_combout ;
wire \F_iw[29]~62_combout ;
wire \F_iw[29]~63_combout ;
wire \D_iw[29]~q ;
wire \E_src1[25]~3_combout ;
wire \F_pc_plus_one[23]~46_combout ;
wire \E_src1[25]~q ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[24]~15_combout ;
wire \F_iw[28]~56_combout ;
wire \F_iw[28]~57_combout ;
wire \D_iw[28]~q ;
wire \E_src1[24]~4_combout ;
wire \F_pc_plus_one[22]~44_combout ;
wire \E_src1[24]~q ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[23]~11_combout ;
wire \F_iw[27]~54_combout ;
wire \F_iw[27]~55_combout ;
wire \D_iw[27]~q ;
wire \E_src1[23]~5_combout ;
wire \F_pc_plus_one[21]~42_combout ;
wire \E_src1[23]~q ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[22]~12_combout ;
wire \F_iw[26]~23_combout ;
wire \F_iw[26]~24_combout ;
wire \D_iw[26]~q ;
wire \E_src1[22]~6_combout ;
wire \F_pc_plus_one[20]~40_combout ;
wire \E_src1[22]~q ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[21]~16_combout ;
wire \F_iw[25]~21_combout ;
wire \F_iw[25]~22_combout ;
wire \D_iw[25]~q ;
wire \E_src1[21]~9_combout ;
wire \F_pc_plus_one[19]~38_combout ;
wire \E_src1[21]~q ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[20]~17_combout ;
wire \F_iw[24]~19_combout ;
wire \F_iw[24]~20_combout ;
wire \D_iw[24]~q ;
wire \E_src1[20]~10_combout ;
wire \F_pc_plus_one[18]~36_combout ;
wire \E_src1[20]~q ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[19]~18_combout ;
wire \F_iw[23]~17_combout ;
wire \F_iw[23]~18_combout ;
wire \D_iw[23]~q ;
wire \E_src1[19]~11_combout ;
wire \F_pc_plus_one[17]~34_combout ;
wire \E_src1[19]~q ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[18]~3_combout ;
wire \F_iw[22]~15_combout ;
wire \F_iw[22]~16_combout ;
wire \D_iw[22]~q ;
wire \E_src1[18]~12_combout ;
wire \F_pc_plus_one[16]~32_combout ;
wire \E_src1[18]~q ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[17]~4_combout ;
wire \F_iw[21]~53_combout ;
wire \D_iw[21]~q ;
wire \E_src1[17]~13_combout ;
wire \F_pc_plus_one[15]~30_combout ;
wire \E_src1[17]~q ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[16]~5_combout ;
wire \F_iw[20]~47_combout ;
wire \D_iw[20]~q ;
wire \E_src1[16]~14_combout ;
wire \F_pc_plus_one[14]~28_combout ;
wire \E_src1[16]~q ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[15]~6_combout ;
wire \F_iw[19]~49_combout ;
wire \F_iw[19]~50_combout ;
wire \D_iw[19]~q ;
wire \E_src1[15]~15_combout ;
wire \F_pc_plus_one[13]~26_combout ;
wire \E_src1[15]~q ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[14]~1_combout ;
wire \F_iw[18]~48_combout ;
wire \F_iw[18]~65_combout ;
wire \D_iw[18]~q ;
wire \E_src1[14]~16_combout ;
wire \F_pc_plus_one[12]~24_combout ;
wire \E_src1[14]~q ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[13]~2_combout ;
wire \F_iw[17]~51_combout ;
wire \F_iw[17]~52_combout ;
wire \F_iw[17]~66_combout ;
wire \D_iw[17]~q ;
wire \E_src1[13]~17_combout ;
wire \F_pc_plus_one[11]~22_combout ;
wire \E_src1[13]~q ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[12]~7_combout ;
wire \E_src1[12]~18_combout ;
wire \F_pc_plus_one[10]~20_combout ;
wire \E_src1[12]~q ;
wire \E_shift_rot_result[12]~q ;
wire \E_shift_rot_result_nxt[11]~8_combout ;
wire \E_src1[11]~19_combout ;
wire \F_pc_plus_one[9]~18_combout ;
wire \E_src1[11]~q ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[10]~9_combout ;
wire \E_src1[10]~20_combout ;
wire \F_pc_plus_one[8]~16_combout ;
wire \E_src1[10]~q ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[9]~10_combout ;
wire \E_src1[9]~21_combout ;
wire \F_pc_plus_one[7]~14_combout ;
wire \E_src1[9]~q ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[8]~13_combout ;
wire \E_src1[8]~22_combout ;
wire \F_pc_plus_one[6]~12_combout ;
wire \E_src1[8]~q ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[7]~0_combout ;
wire \E_shift_rot_result[7]~q ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \Equal0~6_combout ;
wire \D_ctrl_br_cmp~2_combout ;
wire \D_ctrl_br_cmp~5_combout ;
wire \D_ctrl_br_cmp~3_combout ;
wire \D_ctrl_br_cmp~4_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~0_combout ;
wire \R_src2_lo[14]~9_combout ;
wire \E_src2[14]~q ;
wire \Add1~26_combout ;
wire \R_src2_lo[13]~10_combout ;
wire \E_src2[13]~q ;
wire \Add1~27_combout ;
wire \R_src2_lo[12]~11_combout ;
wire \E_src2[12]~q ;
wire \Add1~28_combout ;
wire \R_src2_lo[11]~12_combout ;
wire \E_src2[11]~q ;
wire \Add1~29_combout ;
wire \R_src2_lo[10]~13_combout ;
wire \E_src2[10]~q ;
wire \Add1~30_combout ;
wire \R_src2_lo[9]~14_combout ;
wire \E_src2[9]~q ;
wire \Add1~31_combout ;
wire \R_src2_lo[8]~15_combout ;
wire \E_src2[8]~q ;
wire \Add1~32_combout ;
wire \Add1~25 ;
wire \Add1~34 ;
wire \Add1~36 ;
wire \Add1~38 ;
wire \Add1~40 ;
wire \Add1~42 ;
wire \Add1~44 ;
wire \Add1~45_combout ;
wire \E_logic_result[14]~1_combout ;
wire \W_alu_result[14]~16_combout ;
wire \Add1~43_combout ;
wire \E_logic_result[13]~2_combout ;
wire \W_alu_result[13]~17_combout ;
wire \E_src2[18]~10_combout ;
wire \D_ctrl_unsigned_lo_imm16~3_combout ;
wire \D_ctrl_unsigned_lo_imm16~4_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi~0_combout ;
wire \E_src2[18]~q ;
wire \Add1~47_combout ;
wire \E_src2[17]~11_combout ;
wire \E_src2[17]~q ;
wire \Add1~48_combout ;
wire \E_src2[16]~12_combout ;
wire \E_src2[16]~q ;
wire \Add1~49_combout ;
wire \R_src2_lo[15]~16_combout ;
wire \E_src2[15]~q ;
wire \Add1~50_combout ;
wire \Add1~46 ;
wire \Add1~52 ;
wire \Add1~54 ;
wire \Add1~56 ;
wire \Add1~57_combout ;
wire \E_logic_result[18]~3_combout ;
wire \W_alu_result[18]~12_combout ;
wire \Add1~55_combout ;
wire \E_logic_result[17]~4_combout ;
wire \W_alu_result[17]~13_combout ;
wire \Add1~53_combout ;
wire \E_logic_result[16]~5_combout ;
wire \W_alu_result[16]~14_combout ;
wire \Add1~51_combout ;
wire \E_logic_result[15]~6_combout ;
wire \W_alu_result[15]~15_combout ;
wire \Add1~41_combout ;
wire \E_logic_result[12]~7_combout ;
wire \W_alu_result[12]~18_combout ;
wire \Add1~39_combout ;
wire \E_logic_result[11]~8_combout ;
wire \W_alu_result[11]~19_combout ;
wire \Add1~37_combout ;
wire \E_logic_result[10]~9_combout ;
wire \W_alu_result[10]~20_combout ;
wire \Add1~35_combout ;
wire \E_logic_result[9]~10_combout ;
wire \W_alu_result[9]~21_combout ;
wire \E_src2[23]~5_combout ;
wire \E_src2[23]~q ;
wire \Add1~59_combout ;
wire \E_src2[22]~6_combout ;
wire \E_src2[22]~q ;
wire \Add1~60_combout ;
wire \E_src2[21]~7_combout ;
wire \E_src2[21]~q ;
wire \Add1~61_combout ;
wire \E_src2[20]~8_combout ;
wire \E_src2[20]~q ;
wire \Add1~62_combout ;
wire \E_src2[19]~9_combout ;
wire \E_src2[19]~q ;
wire \Add1~63_combout ;
wire \Add1~58 ;
wire \Add1~65 ;
wire \Add1~67 ;
wire \Add1~69 ;
wire \Add1~71 ;
wire \Add1~72_combout ;
wire \E_logic_result[23]~11_combout ;
wire \W_alu_result[23]~5_combout ;
wire \Add1~70_combout ;
wire \E_logic_result[22]~12_combout ;
wire \W_alu_result[22]~6_combout ;
wire \Add1~33_combout ;
wire \E_logic_result[8]~13_combout ;
wire \W_alu_result[8]~22_combout ;
wire \Add1~22_combout ;
wire \E_logic_result[6]~14_combout ;
wire \W_alu_result[6]~24_combout ;
wire \E_src2[24]~4_combout ;
wire \E_src2[24]~q ;
wire \Add1~74_combout ;
wire \Add1~73 ;
wire \Add1~75_combout ;
wire \E_logic_result[24]~15_combout ;
wire \W_alu_result[24]~4_combout ;
wire \Add1~68_combout ;
wire \E_logic_result[21]~16_combout ;
wire \W_alu_result[21]~9_combout ;
wire \Add1~66_combout ;
wire \E_logic_result[20]~17_combout ;
wire \W_alu_result[20]~10_combout ;
wire \Add1~64_combout ;
wire \E_logic_result[19]~18_combout ;
wire \W_alu_result[19]~11_combout ;
wire \E_src2[28]~0_combout ;
wire \E_src2[28]~q ;
wire \Add1~77_combout ;
wire \E_src2[27]~1_combout ;
wire \E_src2[27]~q ;
wire \Add1~78_combout ;
wire \E_src2[26]~2_combout ;
wire \E_src2[26]~q ;
wire \Add1~79_combout ;
wire \E_src2[25]~3_combout ;
wire \E_src2[25]~q ;
wire \Add1~80_combout ;
wire \Add1~76 ;
wire \Add1~82 ;
wire \Add1~84 ;
wire \Add1~86 ;
wire \Add1~87_combout ;
wire \E_logic_result[28]~19_combout ;
wire \W_alu_result[28]~0_combout ;
wire \Add1~85_combout ;
wire \E_logic_result[27]~20_combout ;
wire \W_alu_result[27]~1_combout ;
wire \Add1~83_combout ;
wire \E_logic_result[26]~21_combout ;
wire \W_alu_result[26]~2_combout ;
wire \Add1~81_combout ;
wire \E_logic_result[25]~22_combout ;
wire \W_alu_result[25]~3_combout ;
wire \Add1~18_combout ;
wire \E_logic_result[4]~23_combout ;
wire \W_alu_result[4]~26_combout ;
wire \Add1~20_combout ;
wire \E_logic_result[5]~24_combout ;
wire \W_alu_result[5]~25_combout ;
wire \Add1~14_combout ;
wire \E_logic_result[2]~25_combout ;
wire \W_alu_result[2]~7_combout ;
wire \Add1~16_combout ;
wire \E_logic_result[3]~26_combout ;
wire \W_alu_result[3]~8_combout ;
wire \d_writedata[24]~0_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \d_writedata[25]~1_combout ;
wire \d_writedata[26]~2_combout ;
wire \d_writedata[27]~3_combout ;
wire \d_writedata[28]~4_combout ;
wire \d_writedata[29]~5_combout ;
wire \d_writedata[30]~6_combout ;
wire \d_writedata[31]~7_combout ;
wire \E_st_stall~combout ;
wire \E_st_data[8]~0_combout ;
wire \E_st_data[9]~1_combout ;
wire \E_st_data[10]~2_combout ;
wire \E_st_data[11]~3_combout ;
wire \E_st_data[12]~4_combout ;
wire \E_st_data[13]~5_combout ;
wire \E_st_data[14]~6_combout ;
wire \E_st_data[15]~7_combout ;
wire \d_writedata[23]~8_combout ;
wire \E_st_data[16]~8_combout ;
wire \E_st_data[17]~9_combout ;
wire \d_read_nxt~0_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \D_ctrl_uncond_cti_non_br~2_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~20_combout ;
wire \R_ctrl_br_uncond~q ;
wire \R_compare_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \R_compare_op[0]~q ;
wire \Equal127~0_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \Equal127~3_combout ;
wire \Equal127~4_combout ;
wire \Equal127~5_combout ;
wire \Equal127~6_combout ;
wire \E_logic_result[0]~27_combout ;
wire \Equal127~7_combout ;
wire \R_src2_hi[15]~1_combout ;
wire \R_src2_hi[15]~2_combout ;
wire \E_src2[31]~q ;
wire \E_logic_result[31]~28_combout ;
wire \E_src2[29]~13_combout ;
wire \E_src2[29]~q ;
wire \E_logic_result[29]~29_combout ;
wire \E_logic_result[1]~30_combout ;
wire \E_src2[30]~14_combout ;
wire \E_src2[30]~q ;
wire \E_logic_result[30]~31_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \E_cmp_result~0_combout ;
wire \E_invert_arith_src_msb~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~q ;
wire \Add1~89_combout ;
wire \E_arith_src1[31]~combout ;
wire \Add1~90_combout ;
wire \Add1~91_combout ;
wire \Add1~88 ;
wire \Add1~93 ;
wire \Add1~95 ;
wire \Add1~97 ;
wire \Add1~98_combout ;
wire \E_cmp_result~1_combout ;
wire \W_cmp_result~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_no_crst_nxt[26]~6_combout ;
wire \F_pc_no_crst_nxt[26]~7_combout ;
wire \F_pc_no_crst_nxt[25]~34_combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \F_pc_no_crst_nxt[25]~8_combout ;
wire \F_pc_no_crst_nxt[24]~9_combout ;
wire \F_pc_no_crst_nxt[23]~10_combout ;
wire \F_pc_no_crst_nxt[22]~35_combout ;
wire \F_pc_no_crst_nxt[22]~11_combout ;
wire \F_pc_no_crst_nxt[21]~12_combout ;
wire \F_pc_no_crst_nxt[20]~13_combout ;
wire \F_pc_no_crst_nxt[19]~14_combout ;
wire \F_pc_no_crst_nxt[18]~15_combout ;
wire \F_pc_no_crst_nxt[17]~16_combout ;
wire \F_pc_no_crst_nxt[16]~17_combout ;
wire \F_pc_no_crst_nxt[15]~18_combout ;
wire \F_pc_no_crst_nxt[14]~19_combout ;
wire \F_pc_no_crst_nxt[13]~20_combout ;
wire \F_pc_no_crst_nxt[12]~21_combout ;
wire \F_pc_no_crst_nxt[11]~22_combout ;
wire \F_pc_no_crst_nxt[10]~23_combout ;
wire \F_pc_no_crst_nxt[9]~36_combout ;
wire \F_pc_no_crst_nxt[9]~24_combout ;
wire \F_pc_no_crst_nxt[8]~25_combout ;
wire \F_pc_no_crst_nxt[7]~26_combout ;
wire \F_pc_no_crst_nxt[5]~27_combout ;
wire \F_pc_no_crst_nxt[6]~28_combout ;
wire \F_pc_no_crst_nxt[4]~29_combout ;
wire \F_pc_no_crst_nxt[1]~30_combout ;
wire \F_pc_no_crst_nxt[3]~31_combout ;
wire \i_read_nxt~0_combout ;
wire \F_pc_no_crst_nxt[2]~32_combout ;
wire \F_pc_no_crst_nxt[0]~33_combout ;
wire \hbreak_enabled~0_combout ;
wire \Add1~10_combout ;
wire \Add1~12_combout ;
wire \E_mem_byte_en[0]~0_combout ;
wire \E_mem_byte_en[1]~1_combout ;
wire \E_mem_byte_en[2]~2_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \E_st_data[18]~10_combout ;
wire \E_st_data[19]~11_combout ;
wire \E_st_data[20]~12_combout ;
wire \E_st_data[21]~13_combout ;
wire \E_st_data[22]~14_combout ;
wire \E_st_data[23]~15_combout ;


usb_system_usb_system_cpu_cpu_nios2_oci the_usb_system_cpu_cpu_nios2_oci(
	.sr_0(sr_0),
	.jtag_break(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.readdata_5(readdata_5),
	.readdata_6(readdata_6),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.resetrequest(debug_reset_request),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr1(WideOr11),
	.local_read(local_read),
	.hbreak_enabled(hbreak_enabled1),
	.mem(mem),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.oci_ienable_6(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[6]~q ),
	.oci_ienable_5(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[5]~q ),
	.oci_single_step_mode(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.readdata_4(readdata_4),
	.r_early_rst(r_early_rst),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_11(readdata_11),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_20(readdata_20),
	.readdata_18(readdata_18),
	.readdata_19(readdata_19),
	.readdata_17(readdata_17),
	.readdata_21(readdata_21),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_31(readdata_31),
	.readdata_30(readdata_30),
	.readdata_29(readdata_29),
	.debugaccess_nxt(src_payload13),
	.writedata_nxt({src_payload43,src_payload44,src_payload45,src_payload42,src_payload41,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload37,src_payload39,src_payload38,src_payload40,src_payload29,src_payload32,src_payload31,src_payload28,
src_payload30,src_payload27,src_payload33,src_payload34,src_payload35,src_payload36,src_payload15,src_payload16,src_payload20,src_payload17,src_payload19,src_payload18,src_payload14}),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_register_bank_b_module usb_system_cpu_cpu_register_bank_b(
	.q_b_0(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_8(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_9(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_10(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_11(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_12(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_15(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_16(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_17(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_18(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_23(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_24(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_28(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_31(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_29(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.D_iw_22(\D_iw[22]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_26(\D_iw[26]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~3_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~4_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~5_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~6_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~8_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~10_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~11_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~12_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~13_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~14_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~15_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~16_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~17_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~18_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~19_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~20_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~21_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~22_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~23_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~24_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~25_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~26_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~27_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~28_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~29_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~30_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~31_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~32_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~33_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~34_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~35_combout ),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_register_bank_a_module usb_system_cpu_cpu_register_bank_a(
	.q_b_7(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_1(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_14(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_18(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_23(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_24(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_28(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_31(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_29(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.D_iw_27(\D_iw[27]~q ),
	.D_iw_28(\D_iw[28]~q ),
	.D_iw_31(\D_iw[31]~q ),
	.D_iw_30(\D_iw[30]~q ),
	.D_iw_29(\D_iw[29]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~3_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~4_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~5_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~6_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~8_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~10_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~11_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~12_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~13_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~14_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~15_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~16_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~17_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~18_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~19_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~20_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~21_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~22_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~23_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~24_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~25_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~26_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~27_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~28_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~29_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~30_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~31_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~32_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~33_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~34_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~35_combout ),
	.clk_clk(clk_clk));

dffeas \W_alu_result[0] (
	.clk(clk_clk),
	.d(\W_alu_result[0]~27_combout ),
	.asdata(\E_shift_rot_result[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

dffeas \W_alu_result[1] (
	.clk(clk_clk),
	.d(\W_alu_result[1]~28_combout ),
	.asdata(\E_shift_rot_result[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

dffeas \av_ld_byte1_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[0]~0_combout ),
	.asdata(\av_ld_byte2_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

dffeas \av_ld_byte1_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[1]~1_combout ),
	.asdata(\av_ld_byte2_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

dffeas \av_ld_byte1_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[2]~2_combout ),
	.asdata(\av_ld_byte2_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

dffeas \av_ld_byte1_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[3]~3_combout ),
	.asdata(\av_ld_byte2_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

dffeas \av_ld_byte1_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[4]~4_combout ),
	.asdata(\av_ld_byte2_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

dffeas \av_ld_byte1_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[5]~5_combout ),
	.asdata(\av_ld_byte2_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

dffeas \av_ld_byte1_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[6]~6_combout ),
	.asdata(\av_ld_byte2_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

dffeas \av_ld_byte1_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[7]~7_combout ),
	.asdata(\av_ld_byte2_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

dffeas \av_ld_byte2_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[0]~0_combout ),
	.asdata(\av_ld_byte3_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

dffeas \av_ld_byte2_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[1]~1_combout ),
	.asdata(\av_ld_byte3_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

cycloneive_lcell_comb \Add1~92 (
	.dataa(\Add1~91_combout ),
	.datab(\E_src1[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~88 ),
	.combout(\Add1~92_combout ),
	.cout(\Add1~93 ));
defparam \Add1~92 .lut_mask = 16'h96EF;
defparam \Add1~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~94 (
	.dataa(\Add1~90_combout ),
	.datab(\E_src1[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~93 ),
	.combout(\Add1~94_combout ),
	.cout(\Add1~95 ));
defparam \Add1~94 .lut_mask = 16'h967F;
defparam \Add1~94 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~96 (
	.dataa(\Add1~89_combout ),
	.datab(\E_arith_src1[31]~combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~95 ),
	.combout(\Add1~96_combout ),
	.cout(\Add1~97 ));
defparam \Add1~96 .lut_mask = 16'h96EF;
defparam \Add1~96 .sum_lutc_input = "cin";

cycloneive_lcell_comb \W_alu_result[0]~27 (
	.dataa(\Add1~10_combout ),
	.datab(\E_logic_result[0]~27_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[0]~27_combout ),
	.cout());
defparam \W_alu_result[0]~27 .lut_mask = 16'hAACC;
defparam \W_alu_result[0]~27 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[2]~4_combout ),
	.asdata(\av_ld_byte3_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

dffeas \av_ld_byte2_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[7]~2_combout ),
	.asdata(\av_ld_byte3_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

dffeas \av_ld_byte2_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[6]~3_combout ),
	.asdata(\av_ld_byte3_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

dffeas \av_ld_byte2_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[5]~7_combout ),
	.asdata(\av_ld_byte3_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

dffeas \av_ld_byte2_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[4]~6_combout ),
	.asdata(\av_ld_byte3_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

dffeas \av_ld_byte2_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[3]~5_combout ),
	.asdata(\av_ld_byte3_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

cycloneive_lcell_comb \W_alu_result[1]~28 (
	.dataa(\Add1~12_combout ),
	.datab(\E_logic_result[1]~30_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[1]~28_combout ),
	.cout());
defparam \W_alu_result[1]~28 .lut_mask = 16'hAACC;
defparam \W_alu_result[1]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[0]~0 (
	.dataa(src_data_8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte1_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[1]~1 (
	.dataa(src_data_9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[1]~1_combout ),
	.cout());
defparam \av_ld_byte1_data[1]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[2]~2 (
	.dataa(src_data_10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[2]~2_combout ),
	.cout());
defparam \av_ld_byte1_data[2]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[3]~3 (
	.dataa(src_data_11),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[3]~3_combout ),
	.cout());
defparam \av_ld_byte1_data[3]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[4]~4 (
	.dataa(src_data_12),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[4]~4_combout ),
	.cout());
defparam \av_ld_byte1_data[4]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[5]~5 (
	.dataa(src_data_13),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[5]~5_combout ),
	.cout());
defparam \av_ld_byte1_data[5]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[6]~6 (
	.dataa(src_data_14),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[6]~6_combout ),
	.cout());
defparam \av_ld_byte1_data[6]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[7]~7 (
	.dataa(src_data_15),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[7]~7_combout ),
	.cout());
defparam \av_ld_byte1_data[7]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[0]~0 (
	.dataa(src_data_16),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte2_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[1]~1 (
	.dataa(src_data_17),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[1]~1_combout ),
	.cout());
defparam \av_ld_byte2_data[1]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[2]~4 (
	.dataa(src_payload7),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[2]~4_combout ),
	.cout());
defparam \av_ld_byte2_data[2]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[7]~2 (
	.dataa(src_payload8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[7]~2_combout ),
	.cout());
defparam \av_ld_byte2_data[7]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[7]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[6]~3 (
	.dataa(src_payload9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[6]~3_combout ),
	.cout());
defparam \av_ld_byte2_data[6]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[6]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[5]~7 (
	.dataa(src_payload10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[5]~7_combout ),
	.cout());
defparam \av_ld_byte2_data[5]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[5]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[4]~6 (
	.dataa(src_payload11),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[4]~6_combout ),
	.cout());
defparam \av_ld_byte2_data[4]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[4]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[3]~5 (
	.dataa(src_payload12),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[3]~5_combout ),
	.cout());
defparam \av_ld_byte2_data[3]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[3]~5 .sum_lutc_input = "datac";

dffeas \W_alu_result[31] (
	.clk(clk_clk),
	.d(\W_alu_result[31]~29_combout ),
	.asdata(\E_shift_rot_result[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(clk_clk),
	.d(\W_alu_result[29]~30_combout ),
	.asdata(\E_shift_rot_result[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(clk_clk),
	.d(\W_alu_result[30]~31_combout ),
	.asdata(\E_shift_rot_result[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

cycloneive_lcell_comb \W_alu_result[31]~29 (
	.dataa(\Add1~96_combout ),
	.datab(\E_logic_result[31]~28_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[31]~29_combout ),
	.cout());
defparam \W_alu_result[31]~29 .lut_mask = 16'hAACC;
defparam \W_alu_result[31]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[29]~30 (
	.dataa(\Add1~92_combout ),
	.datab(\E_logic_result[29]~29_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[29]~30_combout ),
	.cout());
defparam \W_alu_result[29]~30 .lut_mask = 16'hAACC;
defparam \W_alu_result[29]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[30]~31 (
	.dataa(\Add1~94_combout ),
	.datab(\E_logic_result[30]~31_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[30]~31_combout ),
	.cout());
defparam \W_alu_result[30]~31 .lut_mask = 16'hAACC;
defparam \W_alu_result[30]~31 .sum_lutc_input = "datac";

dffeas R_wr_dst_reg(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cycloneive_lcell_comb W_rf_wren(
	.dataa(r_sync_rst),
	.datab(\R_wr_dst_reg~q ),
	.datac(\W_valid~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wren~combout ),
	.cout());
defparam W_rf_wren.lut_mask = 16'hFEFE;
defparam W_rf_wren.sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[0]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~0 (
	.dataa(\R_ctrl_br_cmp~q ),
	.datab(\W_cmp_result~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~0_combout ),
	.cout());
defparam \W_rf_wr_data[0]~0 .lut_mask = 16'hEEEE;
defparam \W_rf_wr_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_control_rd_data[0] (
	.clk(clk_clk),
	.d(\E_control_rd_data[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~1 (
	.dataa(\W_control_rd_data[0]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~1_combout ),
	.cout());
defparam \W_rf_wr_data[0]~1 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[0]~2 (
	.dataa(\av_ld_byte0_data[0]~q ),
	.datab(\W_rf_wr_data[0]~0_combout ),
	.datac(\W_rf_wr_data[0]~1_combout ),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~2_combout ),
	.cout());
defparam \W_rf_wr_data[0]~2 .lut_mask = 16'hFAFC;
defparam \W_rf_wr_data[0]~2 .sum_lutc_input = "datac";

dffeas \R_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

dffeas \av_ld_byte0_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[1]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[1]~3 (
	.dataa(\av_ld_byte0_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[1]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~3_combout ),
	.cout());
defparam \W_rf_wr_data[1]~3 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[1]~3 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[2]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[2]~4 (
	.dataa(\av_ld_byte0_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_2),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[2]~4_combout ),
	.cout());
defparam \W_rf_wr_data[2]~4 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[2]~4 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[3]~5 (
	.dataa(\av_ld_byte0_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_3),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[3]~5_combout ),
	.cout());
defparam \W_rf_wr_data[3]~5 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[3]~5 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[4]~6 (
	.dataa(\av_ld_byte0_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_4),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[4]~6_combout ),
	.cout());
defparam \W_rf_wr_data[4]~6 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[4]~6 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

dffeas \W_control_rd_data[5] (
	.clk(clk_clk),
	.d(\E_control_rd_data[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[5]~q ),
	.prn(vcc));
defparam \W_control_rd_data[5] .is_wysiwyg = "true";
defparam \W_control_rd_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[5]~7 (
	.dataa(\W_control_rd_data[5]~q ),
	.datab(W_alu_result_5),
	.datac(gnd),
	.datad(\R_ctrl_rd_ctl_reg~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[5]~7_combout ),
	.cout());
defparam \W_rf_wr_data[5]~7 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[5]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[5]~8 (
	.dataa(\av_ld_byte0_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_rf_wr_data[5]~7_combout ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[5]~8_combout ),
	.cout());
defparam \W_rf_wr_data[5]~8 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[5]~8 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[6]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

dffeas \W_control_rd_data[6] (
	.clk(clk_clk),
	.d(\E_control_rd_data[6]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[6]~q ),
	.prn(vcc));
defparam \W_control_rd_data[6] .is_wysiwyg = "true";
defparam \W_control_rd_data[6] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[6]~9 (
	.dataa(\W_control_rd_data[6]~q ),
	.datab(W_alu_result_6),
	.datac(gnd),
	.datad(\R_ctrl_rd_ctl_reg~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[6]~9_combout ),
	.cout());
defparam \W_rf_wr_data[6]~9 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[6]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[6]~10 (
	.dataa(\av_ld_byte0_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_rf_wr_data[6]~9_combout ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[6]~10_combout ),
	.cout());
defparam \W_rf_wr_data[6]~10 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[6]~10 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[7]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[4]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[7]~11 (
	.dataa(\av_ld_byte0_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_7),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[7]~11_combout ),
	.cout());
defparam \W_rf_wr_data[7]~11 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[7]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[8]~12 (
	.dataa(\av_ld_byte1_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_8),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[8]~12_combout ),
	.cout());
defparam \W_rf_wr_data[8]~12 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[8]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[9]~13 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_9),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[9]~13_combout ),
	.cout());
defparam \W_rf_wr_data[9]~13 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[9]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[10]~14 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_10),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[10]~14_combout ),
	.cout());
defparam \W_rf_wr_data[10]~14 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[10]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[11]~15 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_11),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[11]~15_combout ),
	.cout());
defparam \W_rf_wr_data[11]~15 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[11]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[12]~16 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_12),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[12]~16_combout ),
	.cout());
defparam \W_rf_wr_data[12]~16 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[12]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[13]~17 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_13),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[13]~17_combout ),
	.cout());
defparam \W_rf_wr_data[13]~17 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[13]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[14]~18 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_14),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[14]~18_combout ),
	.cout());
defparam \W_rf_wr_data[14]~18 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[14]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[15]~19 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_15),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[15]~19_combout ),
	.cout());
defparam \W_rf_wr_data[15]~19 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[15]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[16]~20 (
	.dataa(\av_ld_byte2_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_16),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[16]~20_combout ),
	.cout());
defparam \W_rf_wr_data[16]~20 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[16]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[17]~21 (
	.dataa(\av_ld_byte2_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_17),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[17]~21_combout ),
	.cout());
defparam \W_rf_wr_data[17]~21 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[17]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~0 (
	.dataa(\Equal0~11_combout ),
	.datab(\Equal0~12_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.cout());
defparam \D_wr_dst_reg~0 .lut_mask = 16'hEFFF;
defparam \D_wr_dst_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~1 (
	.dataa(\Equal0~13_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~1_combout ),
	.cout());
defparam \D_wr_dst_reg~1 .lut_mask = 16'hFEFF;
defparam \D_wr_dst_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~14 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\Equal0~14_combout ),
	.cout());
defparam \Equal0~14 .lut_mask = 16'hAFFF;
defparam \Equal0~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 16'hFBFF;
defparam \D_ctrl_implicit_dst_eretaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~1 (
	.dataa(\D_iw[16]~q ),
	.datab(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~1_combout ),
	.cout());
defparam \D_dst_regnum[0]~1 .lut_mask = 16'hEEFF;
defparam \D_dst_regnum[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~2 (
	.dataa(\Equal62~8_combout ),
	.datab(\Equal62~9_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~2_combout ),
	.cout());
defparam \D_dst_regnum[0]~2 .lut_mask = 16'hEFFE;
defparam \D_dst_regnum[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~3 (
	.dataa(\Equal0~14_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\D_dst_regnum[0]~1_combout ),
	.datad(\D_dst_regnum[0]~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~3_combout ),
	.cout());
defparam \D_dst_regnum[0]~3 .lut_mask = 16'hFFFE;
defparam \D_dst_regnum[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~12 (
	.dataa(\D_dst_regnum[0]~3_combout ),
	.datab(\D_dst_regnum[0]~21_combout ),
	.datac(\D_dst_regnum[0]~11_combout ),
	.datad(\D_ctrl_exception~3_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~12_combout ),
	.cout());
defparam \D_dst_regnum[0]~12 .lut_mask = 16'hBFFF;
defparam \D_dst_regnum[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~13 (
	.dataa(\D_dst_regnum[0]~12_combout ),
	.datab(\D_iw[22]~q ),
	.datac(\D_iw[17]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~13_combout ),
	.cout());
defparam \D_dst_regnum[0]~13 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[0]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~14 (
	.dataa(\D_dst_regnum[0]~12_combout ),
	.datab(\D_iw[24]~q ),
	.datac(\D_iw[19]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~14_combout ),
	.cout());
defparam \D_dst_regnum[2]~14 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[2]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[3]~15 (
	.dataa(\D_dst_regnum[0]~12_combout ),
	.datab(\D_iw[25]~q ),
	.datac(\D_iw[20]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~15_combout ),
	.cout());
defparam \D_dst_regnum[3]~15 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[3]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~16 (
	.dataa(\D_dst_regnum[0]~12_combout ),
	.datab(\D_iw[26]~q ),
	.datac(\D_iw[21]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~16_combout ),
	.cout());
defparam \D_dst_regnum[4]~16 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[4]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~18 (
	.dataa(\D_dst_regnum[0]~13_combout ),
	.datab(\D_dst_regnum[2]~14_combout ),
	.datac(\D_dst_regnum[3]~15_combout ),
	.datad(\D_dst_regnum[4]~16_combout ),
	.cin(gnd),
	.combout(\Equal0~18_combout ),
	.cout());
defparam \Equal0~18 .lut_mask = 16'h7FFF;
defparam \Equal0~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~17 (
	.dataa(\D_iw[23]~q ),
	.datab(\D_iw[18]~q ),
	.datac(gnd),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~17_combout ),
	.cout());
defparam \D_dst_regnum[1]~17 .lut_mask = 16'hAACC;
defparam \D_dst_regnum[1]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~18 (
	.dataa(\Equal0~14_combout ),
	.datab(\D_dst_regnum[1]~17_combout ),
	.datac(gnd),
	.datad(\D_dst_regnum[0]~12_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~18_combout ),
	.cout());
defparam \D_dst_regnum[1]~18 .lut_mask = 16'hEEFF;
defparam \D_dst_regnum[1]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~2 (
	.dataa(\D_wr_dst_reg~0_combout ),
	.datab(\D_wr_dst_reg~1_combout ),
	.datac(\Equal0~18_combout ),
	.datad(\D_dst_regnum[1]~18_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~2_combout ),
	.cout());
defparam \D_wr_dst_reg~2 .lut_mask = 16'hFF7F;
defparam \D_wr_dst_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~0 (
	.dataa(\W_alu_result[1]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.cout());
defparam \av_ld_rshift8~0 .lut_mask = 16'hEFFF;
defparam \av_ld_rshift8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~1 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_rshift8~1_combout ),
	.cout());
defparam \av_ld_rshift8~1 .lut_mask = 16'hEEEE;
defparam \av_ld_rshift8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data[4]~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\av_ld_rshift8~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data[4]~0_combout ),
	.cout());
defparam \av_ld_byte0_data[4]~0 .lut_mask = 16'hFF55;
defparam \av_ld_byte0_data[4]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\D_iw[6]~q ),
	.datac(\D_iw[7]~q ),
	.datad(\W_bstatus_reg~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.cout());
defparam \E_control_rd_data[0]~0 .lut_mask = 16'hFFBE;
defparam \E_control_rd_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~1 (
	.dataa(\W_estatus_reg~q ),
	.datab(\D_iw[8]~q ),
	.datac(\D_iw[6]~q ),
	.datad(\E_control_rd_data[0]~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~1_combout ),
	.cout());
defparam \E_control_rd_data[0]~1 .lut_mask = 16'hBFFB;
defparam \E_control_rd_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld_signed~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~1_combout ),
	.cout());
defparam \D_ctrl_ld_signed~1 .lut_mask = 16'hEEEE;
defparam \D_ctrl_ld_signed~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[18]~22 (
	.dataa(\av_ld_byte2_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_18),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[18]~22_combout ),
	.cout());
defparam \W_rf_wr_data[18]~22 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[18]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[23]~23 (
	.dataa(\av_ld_byte2_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_23),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[23]~23_combout ),
	.cout());
defparam \W_rf_wr_data[23]~23 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[23]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[22]~24 (
	.dataa(\av_ld_byte2_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_22),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[22]~24_combout ),
	.cout());
defparam \W_rf_wr_data[22]~24 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[22]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[21]~25 (
	.dataa(\av_ld_byte2_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_21),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[21]~25_combout ),
	.cout());
defparam \W_rf_wr_data[21]~25 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[21]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[20]~26 (
	.dataa(\av_ld_byte2_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_20),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[20]~26_combout ),
	.cout());
defparam \W_rf_wr_data[20]~26 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[20]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[19]~27 (
	.dataa(\av_ld_byte2_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_19),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[19]~27_combout ),
	.cout());
defparam \W_rf_wr_data[19]~27 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[19]~27 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[24]~28 (
	.dataa(\av_ld_byte3_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_24),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[24]~28_combout ),
	.cout());
defparam \W_rf_wr_data[24]~28 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[24]~28 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[28]~29 (
	.dataa(\av_ld_byte3_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_28),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[28]~29_combout ),
	.cout());
defparam \W_rf_wr_data[28]~29 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[28]~29 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[27]~30 (
	.dataa(\av_ld_byte3_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_27),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[27]~30_combout ),
	.cout());
defparam \W_rf_wr_data[27]~30 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[27]~30 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[26]~31 (
	.dataa(\av_ld_byte3_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_26),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[26]~31_combout ),
	.cout());
defparam \W_rf_wr_data[26]~31 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[26]~31 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[25]~32 (
	.dataa(\av_ld_byte3_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_25),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[25]~32_combout ),
	.cout());
defparam \W_rf_wr_data[25]~32 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[25]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~4 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(src_data_2),
	.datac(src_data_21),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~4_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~4 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~5 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(src_data_3),
	.datac(src_data_31),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~5_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~5 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[3]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~6 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(src_data_4),
	.datac(src_data_47),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~6_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~6 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[4]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~7 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(src_data_5),
	.datac(src_data_51),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~7_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~7 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[5]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[5]~2 (
	.dataa(gnd),
	.datab(\D_iw[7]~q ),
	.datac(\D_iw[6]~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[5]~2_combout ),
	.cout());
defparam \E_control_rd_data[5]~2 .lut_mask = 16'hC33C;
defparam \E_control_rd_data[5]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[5]~3 (
	.dataa(\E_control_rd_data[5]~2_combout ),
	.datab(\W_ipending_reg[5]~q ),
	.datac(\W_ienable_reg[5]~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[5]~3_combout ),
	.cout());
defparam \E_control_rd_data[5]~3 .lut_mask = 16'hFAFC;
defparam \E_control_rd_data[5]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~8 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(src_data_6),
	.datac(src_data_61),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~8_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~8 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[6]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[6]~4 (
	.dataa(\E_control_rd_data[5]~2_combout ),
	.datab(\W_ipending_reg[6]~q ),
	.datac(\W_ienable_reg[6]~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[6]~4_combout ),
	.cout());
defparam \E_control_rd_data[6]~4 .lut_mask = 16'hFAFC;
defparam \E_control_rd_data[6]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~9 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(src_data_7),
	.datac(src_data_71),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~9_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~9 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[7]~9 .sum_lutc_input = "datac";

dffeas R_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_ld_signed~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cycloneive_lcell_comb \av_fill_bit~0 (
	.dataa(\R_ctrl_ld_signed~q ),
	.datab(\av_ld_byte1_data[7]~q ),
	.datac(\av_ld_byte0_data[7]~q ),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\av_fill_bit~0_combout ),
	.cout());
defparam \av_fill_bit~0 .lut_mask = 16'hFAFC;
defparam \av_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\D_ctrl_mem16~0_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.cout());
defparam \av_ld_byte1_data_en~0 .lut_mask = 16'hEFFF;
defparam \av_ld_byte1_data_en~0 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

dffeas \av_ld_byte3_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

dffeas \av_ld_byte3_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~0 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_241),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~0_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~0 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~1 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(src_payload6),
	.datac(\av_ld_byte3_data_nxt~0_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~1_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~1 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~2 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_281),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~2_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~2 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~3 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(src_payload6),
	.datac(\av_ld_byte3_data_nxt~2_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~3_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~3 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~4 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_271),
	.datad(av_readdata_pre_27),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~4_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~4 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~5 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~4_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~5_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~6 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_261),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~6_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~6 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~7 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(src_payload6),
	.datac(\av_ld_byte3_data_nxt~6_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~7_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~7 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~8 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_251),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~8_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~8 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~9 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~8_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~9_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~9 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[31]~33 (
	.dataa(\av_ld_byte3_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[31]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[31]~33_combout ),
	.cout());
defparam \W_rf_wr_data[31]~33 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[31]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[29]~34 (
	.dataa(\av_ld_byte3_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[29]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[29]~34_combout ),
	.cout());
defparam \W_rf_wr_data[29]~34 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[29]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[30]~35 (
	.dataa(\av_ld_byte3_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[30]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[30]~35_combout ),
	.cout());
defparam \W_rf_wr_data[30]~35 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[30]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~10 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_311),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~10_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~10 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~11 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~10_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~11_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~11 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~12 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_301),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~12_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~12 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~13 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(src_payload6),
	.datac(\av_ld_byte3_data_nxt~12_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~13_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~13 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~14 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_291),
	.datad(av_readdata_pre_29),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~14_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~14 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~15 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~14_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~15_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~15 .lut_mask = 16'hAACC;
defparam \av_ld_byte3_data_nxt~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~10 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[0]~q ),
	.datad(src_data_0),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~10_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~10 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~11 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[1]~q ),
	.datad(src_data_1),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~11_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~11 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[1]~11 .sum_lutc_input = "datac";

dffeas \W_alu_result[7] (
	.clk(clk_clk),
	.d(\W_alu_result[7]~23_combout ),
	.asdata(\E_shift_rot_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(clk_clk),
	.d(\W_alu_result[14]~16_combout ),
	.asdata(\E_shift_rot_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(clk_clk),
	.d(\W_alu_result[13]~17_combout ),
	.asdata(\E_shift_rot_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(clk_clk),
	.d(\W_alu_result[18]~12_combout ),
	.asdata(\E_shift_rot_result[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_18),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(clk_clk),
	.d(\W_alu_result[17]~13_combout ),
	.asdata(\E_shift_rot_result[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_17),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(clk_clk),
	.d(\W_alu_result[16]~14_combout ),
	.asdata(\E_shift_rot_result[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_16),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(clk_clk),
	.d(\W_alu_result[15]~15_combout ),
	.asdata(\E_shift_rot_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[12] (
	.clk(clk_clk),
	.d(\W_alu_result[12]~18_combout ),
	.asdata(\E_shift_rot_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(clk_clk),
	.d(\W_alu_result[11]~19_combout ),
	.asdata(\E_shift_rot_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(clk_clk),
	.d(\W_alu_result[10]~20_combout ),
	.asdata(\E_shift_rot_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(clk_clk),
	.d(\W_alu_result[9]~21_combout ),
	.asdata(\E_shift_rot_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(clk_clk),
	.d(\W_alu_result[23]~5_combout ),
	.asdata(\E_shift_rot_result[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_23),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(clk_clk),
	.d(\W_alu_result[22]~6_combout ),
	.asdata(\E_shift_rot_result[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_22),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(clk_clk),
	.d(\W_alu_result[8]~22_combout ),
	.asdata(\E_shift_rot_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[6] (
	.clk(clk_clk),
	.d(\W_alu_result[6]~24_combout ),
	.asdata(\E_shift_rot_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(clk_clk),
	.d(\W_alu_result[24]~4_combout ),
	.asdata(\E_shift_rot_result[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_24),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(clk_clk),
	.d(\W_alu_result[21]~9_combout ),
	.asdata(\E_shift_rot_result[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_21),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(clk_clk),
	.d(\W_alu_result[20]~10_combout ),
	.asdata(\E_shift_rot_result[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_20),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(clk_clk),
	.d(\W_alu_result[19]~11_combout ),
	.asdata(\E_shift_rot_result[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_19),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \W_alu_result[28] (
	.clk(clk_clk),
	.d(\W_alu_result[28]~0_combout ),
	.asdata(\E_shift_rot_result[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_28),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \W_alu_result[27] (
	.clk(clk_clk),
	.d(\W_alu_result[27]~1_combout ),
	.asdata(\E_shift_rot_result[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_27),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(clk_clk),
	.d(\W_alu_result[26]~2_combout ),
	.asdata(\E_shift_rot_result[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_26),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(clk_clk),
	.d(\W_alu_result[25]~3_combout ),
	.asdata(\E_shift_rot_result[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_25),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \W_alu_result[4] (
	.clk(clk_clk),
	.d(\W_alu_result[4]~26_combout ),
	.asdata(\E_shift_rot_result[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(clk_clk),
	.d(\W_alu_result[5]~25_combout ),
	.asdata(\E_shift_rot_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(clk_clk),
	.d(\W_alu_result[2]~7_combout ),
	.asdata(\E_shift_rot_result[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(clk_clk),
	.d(\W_alu_result[3]~8_combout ),
	.asdata(\E_shift_rot_result[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\d_writedata[24]~0_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\d_writedata[25]~1_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\d_writedata[26]~2_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\d_writedata[27]~3_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\d_writedata[28]~4_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\d_writedata[29]~5_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\d_writedata[30]~6_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\d_writedata[31]~7_combout ),
	.asdata(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\E_st_data[8]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\E_st_data[9]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\E_st_data[10]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\E_st_data[11]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\E_st_data[12]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\E_st_data[13]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\E_st_data[14]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\E_st_data[15]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\E_st_data[16]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\E_st_data[17]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

cycloneive_lcell_comb \av_ld_getting_data~6 (
	.dataa(WideOr1),
	.datab(\av_ld_getting_data~2_combout ),
	.datac(\av_ld_getting_data~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_ld_getting_data),
	.cout());
defparam \av_ld_getting_data~6 .lut_mask = 16'hFEFE;
defparam \av_ld_getting_data~6 .sum_lutc_input = "datac";

dffeas \F_pc[26] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[26]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_26),
	.prn(vcc));
defparam \F_pc[26] .is_wysiwyg = "true";
defparam \F_pc[26] .power_up = "low";

dffeas \F_pc[25] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[25]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_25),
	.prn(vcc));
defparam \F_pc[25] .is_wysiwyg = "true";
defparam \F_pc[25] .power_up = "low";

dffeas \F_pc[24] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[24]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_24),
	.prn(vcc));
defparam \F_pc[24] .is_wysiwyg = "true";
defparam \F_pc[24] .power_up = "low";

dffeas \F_pc[23] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[23]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_23),
	.prn(vcc));
defparam \F_pc[23] .is_wysiwyg = "true";
defparam \F_pc[23] .power_up = "low";

dffeas \F_pc[22] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[22]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_22),
	.prn(vcc));
defparam \F_pc[22] .is_wysiwyg = "true";
defparam \F_pc[22] .power_up = "low";

dffeas \F_pc[21] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[21]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_21),
	.prn(vcc));
defparam \F_pc[21] .is_wysiwyg = "true";
defparam \F_pc[21] .power_up = "low";

dffeas \F_pc[20] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[20]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_20),
	.prn(vcc));
defparam \F_pc[20] .is_wysiwyg = "true";
defparam \F_pc[20] .power_up = "low";

dffeas \F_pc[19] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[19]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_19),
	.prn(vcc));
defparam \F_pc[19] .is_wysiwyg = "true";
defparam \F_pc[19] .power_up = "low";

dffeas \F_pc[18] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[18]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_18),
	.prn(vcc));
defparam \F_pc[18] .is_wysiwyg = "true";
defparam \F_pc[18] .power_up = "low";

dffeas \F_pc[17] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[17]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_17),
	.prn(vcc));
defparam \F_pc[17] .is_wysiwyg = "true";
defparam \F_pc[17] .power_up = "low";

dffeas \F_pc[16] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[16]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_16),
	.prn(vcc));
defparam \F_pc[16] .is_wysiwyg = "true";
defparam \F_pc[16] .power_up = "low";

dffeas \F_pc[15] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[15]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_15),
	.prn(vcc));
defparam \F_pc[15] .is_wysiwyg = "true";
defparam \F_pc[15] .power_up = "low";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[14]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_14),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[13]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[12]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[11]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[10]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[9]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[8]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[7]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[5]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[6]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[4]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[1]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[3]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[2]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[0]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\E_st_data[18]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\E_st_data[19]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\E_st_data[20]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\E_st_data[21]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\E_st_data[22]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\E_st_data[23]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

cycloneive_lcell_comb \F_valid~0 (
	.dataa(WideOr12),
	.datab(av_readdatavalid),
	.datac(av_readdatavalid1),
	.datad(i_read1),
	.cin(gnd),
	.combout(\F_valid~0_combout ),
	.cout());
defparam \F_valid~0 .lut_mask = 16'hFEFF;
defparam \F_valid~0 .sum_lutc_input = "datac";

dffeas D_valid(
	.clk(clk_clk),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(clk_clk),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

cycloneive_lcell_comb \F_iw[11]~25 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_11),
	.datad(av_readdata_pre_111),
	.cin(gnd),
	.combout(\F_iw[11]~25_combout ),
	.cout());
defparam \F_iw[11]~25 .lut_mask = 16'hFFFE;
defparam \F_iw[11]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~37 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\F_iw[10]~37_combout ),
	.cout());
defparam \F_iw[10]~37 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~38 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[10]~37_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_10),
	.cin(gnd),
	.combout(\F_iw[10]~38_combout ),
	.cout());
defparam \F_iw[10]~38 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~38 .sum_lutc_input = "datac";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cycloneive_lcell_comb \F_iw[4]~13 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_4),
	.datad(av_readdata_pre_4),
	.cin(gnd),
	.combout(\F_iw[4]~13_combout ),
	.cout());
defparam \F_iw[4]~13 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[4]~14 (
	.dataa(\F_iw[4]~13_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[4]~14_combout ),
	.cout());
defparam \F_iw[4]~14 .lut_mask = 16'hFEFF;
defparam \F_iw[4]~14 .sum_lutc_input = "datac";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cycloneive_lcell_comb \F_iw[1]~8 (
	.dataa(src_payload),
	.datab(out_valid2),
	.datac(out_data_buffer_1),
	.datad(av_readdata_pre_1),
	.cin(gnd),
	.combout(\F_iw[1]~8_combout ),
	.cout());
defparam \F_iw[1]~8 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[1]~9 (
	.dataa(\F_iw[1]~8_combout ),
	.datab(src1_valid),
	.datac(av_readdata_pre_11),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[1]~9_combout ),
	.cout());
defparam \F_iw[1]~9 .lut_mask = 16'hFEFF;
defparam \F_iw[1]~9 .sum_lutc_input = "datac";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cycloneive_lcell_comb \F_iw[0]~6 (
	.dataa(src_payload),
	.datab(out_valid2),
	.datac(out_data_buffer_0),
	.datad(av_readdata_pre_0),
	.cin(gnd),
	.combout(\F_iw[0]~6_combout ),
	.cout());
defparam \F_iw[0]~6 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~7 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[0]~6_combout ),
	.datac(src1_valid),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(\F_iw[0]~7_combout ),
	.cout());
defparam \F_iw[0]~7 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~7 .sum_lutc_input = "datac";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cycloneive_lcell_comb \F_iw[3]~12 (
	.dataa(src_payload2),
	.datab(src1_valid),
	.datac(av_readdata_pre_3),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[3]~12_combout ),
	.cout());
defparam \F_iw[3]~12 .lut_mask = 16'hFEFF;
defparam \F_iw[3]~12 .sum_lutc_input = "datac";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cycloneive_lcell_comb \F_iw[2]~10 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_2),
	.datad(av_readdata_pre_2),
	.cin(gnd),
	.combout(\F_iw[2]~10_combout ),
	.cout());
defparam \F_iw[2]~10 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~11 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[2]~10_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[2]~11_combout ),
	.cout());
defparam \F_iw[2]~11 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~11 .sum_lutc_input = "datac";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFBFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~32 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_5),
	.datad(av_readdata_pre_5),
	.cin(gnd),
	.combout(\F_iw[5]~32_combout ),
	.cout());
defparam \F_iw[5]~32 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~33 (
	.dataa(\F_iw[5]~32_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[5]~33_combout ),
	.cout());
defparam \F_iw[5]~33 .lut_mask = 16'hFEFF;
defparam \F_iw[5]~33 .sum_lutc_input = "datac";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cycloneive_lcell_comb \Equal0~7 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~2_combout ),
	.datac(\D_iw[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'hFEFE;
defparam \Equal0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~35 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_15),
	.datad(av_readdata_pre_15),
	.cin(gnd),
	.combout(\F_iw[15]~35_combout ),
	.cout());
defparam \F_iw[15]~35 .lut_mask = 16'hFFFE;
defparam \F_iw[15]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~36 (
	.dataa(\F_iw[15]~35_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[15]~36_combout ),
	.cout());
defparam \F_iw[15]~36 .lut_mask = 16'hFEFF;
defparam \F_iw[15]~36 .sum_lutc_input = "datac";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~36_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

dffeas E_new_inst(
	.clk(clk_clk),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

cycloneive_lcell_comb \D_ctrl_st~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.cout());
defparam \D_ctrl_st~0 .lut_mask = 16'hBFFF;
defparam \D_ctrl_st~0 .sum_lutc_input = "datac";

dffeas R_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cycloneive_lcell_comb \W_valid~3 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\E_valid_from_R~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_valid~3_combout ),
	.cout());
defparam \W_valid~3 .lut_mask = 16'hF7F7;
defparam \W_valid~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_valid~2 (
	.dataa(\E_stall~4_combout ),
	.datab(d_write1),
	.datac(av_waitrequest),
	.datad(\W_valid~3_combout ),
	.cin(gnd),
	.combout(\W_valid~2_combout ),
	.cout());
defparam \W_valid~2 .lut_mask = 16'hFF7F;
defparam \W_valid~2 .sum_lutc_input = "datac";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cycloneive_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(\hbreak_pending~q ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.cout());
defparam \hbreak_pending_nxt~0 .lut_mask = 16'hEEFF;
defparam \hbreak_pending_nxt~0 .sum_lutc_input = "datac";

dffeas hbreak_pending(
	.clk(clk_clk),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cycloneive_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datab(hbreak_enabled1),
	.datac(\wait_for_one_post_bret_inst~q ),
	.datad(\F_valid~0_combout ),
	.cin(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.cout());
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 16'hFEFF;
defparam \wait_for_one_post_bret_inst~0 .sum_lutc_input = "datac";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cycloneive_lcell_comb \hbreak_req~0 (
	.dataa(\W_valid~q ),
	.datab(\hbreak_pending~q ),
	.datac(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.datad(\wait_for_one_post_bret_inst~q ),
	.cin(gnd),
	.combout(\hbreak_req~0_combout ),
	.cout());
defparam \hbreak_req~0 .lut_mask = 16'hFEFF;
defparam \hbreak_req~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~34 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_14),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\F_iw[14]~34_combout ),
	.cout());
defparam \F_iw[14]~34 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~64 (
	.dataa(\D_iw[5]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[14]~34_combout ),
	.cin(gnd),
	.combout(\F_iw[14]~64_combout ),
	.cout());
defparam \F_iw[14]~64 .lut_mask = 16'hFFDF;
defparam \F_iw[14]~64 .sum_lutc_input = "datac";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cycloneive_lcell_comb \D_op_opx_rsv63~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_op_opx_rsv63~0_combout ),
	.cout());
defparam \D_op_opx_rsv63~0 .lut_mask = 16'hEEEE;
defparam \D_op_opx_rsv63~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~27 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_13),
	.datad(av_readdata_pre_13),
	.cin(gnd),
	.combout(\F_iw[13]~27_combout ),
	.cout());
defparam \F_iw[13]~27 .lut_mask = 16'hFFFE;
defparam \F_iw[13]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~28 (
	.dataa(\F_iw[13]~27_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[13]~28_combout ),
	.cout());
defparam \F_iw[13]~28 .lut_mask = 16'hFEFF;
defparam \F_iw[13]~28 .sum_lutc_input = "datac";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

cycloneive_lcell_comb \F_iw[16]~29 (
	.dataa(src_payload3),
	.datab(src1_valid),
	.datac(av_readdata_pre_16),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[16]~29_combout ),
	.cout());
defparam \F_iw[16]~29 .lut_mask = 16'hFEFF;
defparam \F_iw[16]~29 .sum_lutc_input = "datac";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cycloneive_lcell_comb \F_iw[12]~30 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_12),
	.cin(gnd),
	.combout(\F_iw[12]~30_combout ),
	.cout());
defparam \F_iw[12]~30 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[12]~31 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[12]~30_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_12),
	.cin(gnd),
	.combout(\F_iw[12]~31_combout ),
	.cout());
defparam \F_iw[12]~31 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~31 .sum_lutc_input = "datac";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cycloneive_lcell_comb \Equal62~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~4_combout ),
	.cout());
defparam \Equal62~4 .lut_mask = 16'hFF7F;
defparam \Equal62~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~5 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~5_combout ),
	.cout());
defparam \Equal62~5 .lut_mask = 16'hFFF7;
defparam \Equal62~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~6 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~6_combout ),
	.cout());
defparam \Equal62~6 .lut_mask = 16'hFFFB;
defparam \Equal62~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~5_combout ),
	.datad(\Equal62~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~7 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~7_combout ),
	.cout());
defparam \Equal62~7 .lut_mask = 16'hFFBF;
defparam \Equal62~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(\Equal62~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_shift_rot~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(\D_iw[12]~q ),
	.datab(gnd),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.cout());
defparam \D_ctrl_shift_logical~0 .lut_mask = 16'hAFFF;
defparam \D_ctrl_shift_logical~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.cout());
defparam \D_ctrl_shift_rot~2 .lut_mask = 16'hACFF;
defparam \D_ctrl_shift_rot~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~3 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_shift_rot~0_combout ),
	.datac(\D_ctrl_shift_rot~1_combout ),
	.datad(\D_ctrl_shift_rot~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~3_combout ),
	.cout());
defparam \D_ctrl_shift_rot~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~3 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[0]~5 (
	.dataa(\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\E_shift_rot_cnt[0]~5_combout ),
	.cout(\E_shift_rot_cnt[0]~6 ));
defparam \E_shift_rot_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \E_shift_rot_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~0 .lut_mask = 16'hFFF7;
defparam \D_ctrl_hi_imm16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\D_ctrl_hi_imm16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~1_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~1 .lut_mask = 16'hFEFE;
defparam \D_ctrl_hi_imm16~1 .sum_lutc_input = "datac";

dffeas R_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_hi_imm16~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cycloneive_lcell_comb \Equal0~12 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~12_combout ),
	.cout());
defparam \Equal0~12 .lut_mask = 16'hDFFF;
defparam \Equal0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[0]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~14_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~14 .lut_mask = 16'hF6FF;
defparam \D_ctrl_alu_force_xor~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~17 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~17_combout ),
	.cout());
defparam \Equal0~17 .lut_mask = 16'hFFFE;
defparam \Equal0~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~11 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~11_combout ),
	.cout());
defparam \Equal0~11 .lut_mask = 16'hFFFD;
defparam \Equal0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~2 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_ctrl_alu_force_xor~14_combout ),
	.datac(\Equal0~17_combout ),
	.datad(\Equal0~11_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~2_combout ),
	.cout());
defparam \D_ctrl_exception~2 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~14 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~14_combout ),
	.cout());
defparam \Equal62~14 .lut_mask = 16'hFEFF;
defparam \Equal62~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~9 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~9_combout ),
	.cout());
defparam \Equal62~9 .lut_mask = 16'hFDFF;
defparam \Equal62~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~14_combout ),
	.datac(\Equal62~9_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~13 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~13_combout ),
	.cout());
defparam \Equal62~13 .lut_mask = 16'hEFFF;
defparam \Equal62~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal62~13_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~16 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~16_combout ),
	.cout());
defparam \Equal0~16 .lut_mask = 16'hBFFF;
defparam \Equal0~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~16_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 16'hFFDE;
defparam \D_ctrl_force_src2_zero~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~3 (
	.dataa(\D_ctrl_exception~2_combout ),
	.datab(\D_ctrl_force_src2_zero~1_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_force_src2_zero~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~3_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~3 .lut_mask = 16'hFFFD;
defparam \D_ctrl_force_src2_zero~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hEEEE;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv00~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv00~0_combout ),
	.cout());
defparam \D_op_opx_rsv00~0 .lut_mask = 16'hEFFF;
defparam \D_op_opx_rsv00~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~2_combout ),
	.cout());
defparam \Equal62~2 .lut_mask = 16'hFBFF;
defparam \Equal62~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~20 (
	.dataa(\Equal62~0_combout ),
	.datab(\Equal62~2_combout ),
	.datac(\Equal62~6_combout ),
	.datad(\Equal62~5_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~20_combout ),
	.cout());
defparam \D_dst_regnum[0]~20 .lut_mask = 16'h7FFF;
defparam \D_dst_regnum[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~10_combout ),
	.cout());
defparam \Equal62~10 .lut_mask = 16'hBFFF;
defparam \Equal62~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~11 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~11_combout ),
	.cout());
defparam \Equal62~11 .lut_mask = 16'hDFFF;
defparam \Equal62~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv17~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv17~0_combout ),
	.cout());
defparam \D_op_opx_rsv17~0 .lut_mask = 16'hFEFF;
defparam \D_op_opx_rsv17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~5 (
	.dataa(gnd),
	.datab(\Equal62~10_combout ),
	.datac(\Equal62~11_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~5_combout ),
	.cout());
defparam \D_dst_regnum[0]~5 .lut_mask = 16'h3FFF;
defparam \D_dst_regnum[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~8 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~8_combout ),
	.cout());
defparam \Equal62~8 .lut_mask = 16'hFFEF;
defparam \Equal62~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_cmpge~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_cmpge~0_combout ),
	.cout());
defparam \D_op_cmpge~0 .lut_mask = 16'hFEFF;
defparam \D_op_cmpge~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~4 (
	.dataa(gnd),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~8_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~4_combout ),
	.cout());
defparam \D_dst_regnum[0]~4 .lut_mask = 16'h3FFF;
defparam \D_dst_regnum[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~21 (
	.dataa(\D_op_opx_rsv00~0_combout ),
	.datab(\D_dst_regnum[0]~20_combout ),
	.datac(\D_dst_regnum[0]~5_combout ),
	.datad(\D_dst_regnum[0]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~21_combout ),
	.cout());
defparam \D_dst_regnum[0]~21 .lut_mask = 16'hFFFD;
defparam \D_dst_regnum[0]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~15 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~15_combout ),
	.cout());
defparam \Equal0~15 .lut_mask = 16'hFDFF;
defparam \Equal0~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~6 (
	.dataa(\Equal62~5_combout ),
	.datab(\Equal62~6_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~6_combout ),
	.cout());
defparam \D_dst_regnum[0]~6 .lut_mask = 16'h7FFF;
defparam \D_dst_regnum[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~12 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~12_combout ),
	.cout());
defparam \Equal62~12 .lut_mask = 16'hFFFE;
defparam \Equal62~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~7 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~7_combout ),
	.cout());
defparam \D_dst_regnum[0]~7 .lut_mask = 16'h7F7F;
defparam \D_dst_regnum[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~1_combout ),
	.cout());
defparam \Equal62~1 .lut_mask = 16'hF7FF;
defparam \Equal62~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~3 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~3_combout ),
	.cout());
defparam \Equal62~3 .lut_mask = 16'hFFFD;
defparam \Equal62~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~8 (
	.dataa(\Equal62~1_combout ),
	.datab(\Equal62~10_combout ),
	.datac(\Equal62~3_combout ),
	.datad(\Equal62~9_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~8_combout ),
	.cout());
defparam \D_dst_regnum[0]~8 .lut_mask = 16'h7FFF;
defparam \D_dst_regnum[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~9 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_op_opx_rsv63~0_combout ),
	.datac(\D_dst_regnum[0]~7_combout ),
	.datad(\D_dst_regnum[0]~8_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~9_combout ),
	.cout());
defparam \D_dst_regnum[0]~9 .lut_mask = 16'hFFF7;
defparam \D_dst_regnum[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~10 (
	.dataa(\D_op_opx_rsv17~0_combout ),
	.datab(\Equal62~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~10_combout ),
	.cout());
defparam \D_dst_regnum[0]~10 .lut_mask = 16'h7777;
defparam \D_dst_regnum[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~11 (
	.dataa(\Equal0~15_combout ),
	.datab(\D_dst_regnum[0]~6_combout ),
	.datac(\D_dst_regnum[0]~9_combout ),
	.datad(\D_dst_regnum[0]~10_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~11_combout ),
	.cout());
defparam \D_dst_regnum[0]~11 .lut_mask = 16'hFFFD;
defparam \D_dst_regnum[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'h7FFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~0 .lut_mask = 16'h0FFF;
defparam \D_ctrl_jmp_direct~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~11_combout ),
	.datac(\Equal62~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.cout());
defparam \D_ctrl_retaddr~0 .lut_mask = 16'hFEFE;
defparam \D_ctrl_retaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(\Equal62~9_combout ),
	.datab(\Equal62~14_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.cout());
defparam \D_ctrl_retaddr~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_retaddr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_retaddr~0_combout ),
	.datad(\D_ctrl_retaddr~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.cout());
defparam \D_ctrl_retaddr~2 .lut_mask = 16'hFFFE;
defparam \D_ctrl_retaddr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~4 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~16_combout ),
	.datac(\D_ctrl_jmp_direct~0_combout ),
	.datad(\D_ctrl_retaddr~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~4_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~4 .lut_mask = 16'h7FFF;
defparam \D_ctrl_force_src2_zero~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~19 (
	.dataa(\Equal0~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\Equal0~19_combout ),
	.cout());
defparam \Equal0~19 .lut_mask = 16'hAAFF;
defparam \Equal0~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~5 (
	.dataa(\D_dst_regnum[0]~21_combout ),
	.datab(\D_dst_regnum[0]~11_combout ),
	.datac(\D_ctrl_force_src2_zero~4_combout ),
	.datad(\Equal0~19_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~5_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~5 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(\D_iw[15]~q ),
	.datab(gnd),
	.datac(\Equal0~7_combout ),
	.datad(\Equal62~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 16'hAFFF;
defparam \D_ctrl_uncond_cti_non_br~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~6 (
	.dataa(\Equal0~12_combout ),
	.datab(\D_ctrl_force_src2_zero~3_combout ),
	.datac(\D_ctrl_force_src2_zero~5_combout ),
	.datad(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~6_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~6 .lut_mask = 16'hEFFF;
defparam \D_ctrl_force_src2_zero~6 .sum_lutc_input = "datac";

dffeas R_ctrl_force_src2_zero(
	.clk(clk_clk),
	.d(\D_ctrl_force_src2_zero~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

cycloneive_lcell_comb \R_src2_lo[2]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\R_ctrl_hi_imm16~q ),
	.datad(\R_ctrl_force_src2_zero~q ),
	.cin(gnd),
	.combout(\R_src2_lo[2]~3_combout ),
	.cout());
defparam \R_src2_lo[2]~3 .lut_mask = 16'h0FFF;
defparam \R_src2_lo[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~45 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_6),
	.datad(av_readdata_pre_6),
	.cin(gnd),
	.combout(\F_iw[6]~45_combout ),
	.cout());
defparam \F_iw[6]~45 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~46 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[6]~45_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[6]~46_combout ),
	.cout());
defparam \F_iw[6]~46 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~46 .sum_lutc_input = "datac";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cycloneive_lcell_comb \D_dst_regnum[0]~0 (
	.dataa(\D_iw[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~0_combout ),
	.cout());
defparam \D_dst_regnum[0]~0 .lut_mask = 16'hAAFF;
defparam \D_dst_regnum[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~2 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~4_combout ),
	.datad(\D_dst_regnum[0]~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_unsigned_lo_imm16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~5 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~2_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_unsigned_lo_imm16~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~0 .lut_mask = 16'h6996;
defparam \D_ctrl_b_is_dst~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~1_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~1 .lut_mask = 16'hFBFE;
defparam \D_ctrl_b_is_dst~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~2 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_ctrl_b_is_dst~0_combout ),
	.datad(\D_ctrl_b_is_dst~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~2_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~2 .lut_mask = 16'h96FF;
defparam \D_ctrl_b_is_dst~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~13 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~13_combout ),
	.cout());
defparam \Equal0~13 .lut_mask = 16'hFFDF;
defparam \Equal0~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~0 (
	.dataa(\D_ctrl_b_is_dst~2_combout ),
	.datab(\Equal0~13_combout ),
	.datac(\Equal0~11_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.cout());
defparam \R_src2_use_imm~0 .lut_mask = 16'hFEFF;
defparam \R_src2_use_imm~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.cout());
defparam \R_ctrl_br_nxt~0 .lut_mask = 16'hFFFE;
defparam \R_ctrl_br_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~1 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~1_combout ),
	.cout());
defparam \R_ctrl_br_nxt~1 .lut_mask = 16'hEEFF;
defparam \R_ctrl_br_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~1 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\R_src2_use_imm~0_combout ),
	.datac(\R_valid~q ),
	.datad(\R_ctrl_br_nxt~1_combout ),
	.cin(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.cout());
defparam \R_src2_use_imm~1 .lut_mask = 16'hFFFE;
defparam \R_src2_use_imm~1 .sum_lutc_input = "datac";

dffeas R_src2_use_imm(
	.clk(clk_clk),
	.d(\R_src2_use_imm~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 16'hBBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 16'hEFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .sum_lutc_input = "datac";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cycloneive_lcell_comb \E_src2[3]~16 (
	.dataa(\R_src2_use_imm~q ),
	.datab(\R_ctrl_src_imm5_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[3]~16_combout ),
	.cout());
defparam \E_src2[3]~16 .lut_mask = 16'hEEEE;
defparam \E_src2[3]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[0]~8 (
	.dataa(\R_src2_lo[2]~3_combout ),
	.datab(\D_iw[6]~q ),
	.datac(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\E_src2[3]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[0]~8_combout ),
	.cout());
defparam \R_src2_lo[0]~8 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[0]~8 .sum_lutc_input = "datac";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\R_src2_lo[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

dffeas \E_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[0]~5_combout ),
	.asdata(\E_src2[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[1]~7 (
	.dataa(\E_shift_rot_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[0]~6 ),
	.combout(\E_shift_rot_cnt[1]~7_combout ),
	.cout(\E_shift_rot_cnt[1]~8 ));
defparam \E_shift_rot_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[7]~43 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_7),
	.datad(av_readdata_pre_7),
	.cin(gnd),
	.combout(\F_iw[7]~43_combout ),
	.cout());
defparam \F_iw[7]~43 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~44 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[7]~43_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[7]~44_combout ),
	.cout());
defparam \F_iw[7]~44 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~44 .sum_lutc_input = "datac";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[1]~7 (
	.dataa(\R_src2_lo[2]~3_combout ),
	.datab(\D_iw[7]~q ),
	.datac(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\E_src2[3]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[1]~7_combout ),
	.cout());
defparam \R_src2_lo[1]~7 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[1]~7 .sum_lutc_input = "datac";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\R_src2_lo[1]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[1]~7_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[2]~9 (
	.dataa(\E_shift_rot_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[1]~8 ),
	.combout(\E_shift_rot_cnt[2]~9_combout ),
	.cout(\E_shift_rot_cnt[2]~10 ));
defparam \E_shift_rot_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \E_shift_rot_cnt[2]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[8]~41 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_8),
	.datad(av_readdata_pre_8),
	.cin(gnd),
	.combout(\F_iw[8]~41_combout ),
	.cout());
defparam \F_iw[8]~41 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~42 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[8]~41_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[8]~42_combout ),
	.cout());
defparam \F_iw[8]~42 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~42 .sum_lutc_input = "datac";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[2]~6 (
	.dataa(\R_src2_lo[2]~3_combout ),
	.datab(\D_iw[8]~q ),
	.datac(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datad(\E_src2[3]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[2]~6_combout ),
	.cout());
defparam \R_src2_lo[2]~6 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[2]~6 .sum_lutc_input = "datac";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\R_src2_lo[2]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[2]~9_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cycloneive_lcell_comb \E_stall~0 (
	.dataa(\E_new_inst~q ),
	.datab(\E_shift_rot_cnt[0]~q ),
	.datac(\E_shift_rot_cnt[1]~q ),
	.datad(\E_shift_rot_cnt[2]~q ),
	.cin(gnd),
	.combout(\E_stall~0_combout ),
	.cout());
defparam \E_stall~0 .lut_mask = 16'hFFFE;
defparam \E_stall~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_cnt[3]~11 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[2]~10 ),
	.combout(\E_shift_rot_cnt[3]~11_combout ),
	.cout(\E_shift_rot_cnt[3]~12 ));
defparam \E_shift_rot_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[3]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[9]~39 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_9),
	.datad(av_readdata_pre_9),
	.cin(gnd),
	.combout(\F_iw[9]~39_combout ),
	.cout());
defparam \F_iw[9]~39 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[9]~40 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[9]~39_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[9]~40_combout ),
	.cout());
defparam \F_iw[9]~40 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~40 .sum_lutc_input = "datac";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[3]~5 (
	.dataa(\R_src2_lo[2]~3_combout ),
	.datab(\D_iw[9]~q ),
	.datac(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datad(\E_src2[3]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[3]~5_combout ),
	.cout());
defparam \R_src2_lo[3]~5 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[3]~5 .sum_lutc_input = "datac";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\R_src2_lo[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[3]~11_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[4]~13 (
	.dataa(\E_shift_rot_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\E_shift_rot_cnt[3]~12 ),
	.combout(\E_shift_rot_cnt[4]~13_combout ),
	.cout());
defparam \E_shift_rot_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \E_shift_rot_cnt[4]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \R_src2_lo[4]~4 (
	.dataa(\R_src2_lo[2]~3_combout ),
	.datab(\D_iw[10]~q ),
	.datac(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datad(\E_src2[3]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~4_combout ),
	.cout());
defparam \R_src2_lo[4]~4 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[4]~4 .sum_lutc_input = "datac";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\R_src2_lo[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[4]~13_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cycloneive_lcell_comb \E_stall~1 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(\E_shift_rot_cnt[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_stall~1_combout ),
	.cout());
defparam \E_stall~1 .lut_mask = 16'hEEEE;
defparam \E_stall~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~2 (
	.dataa(\R_ctrl_shift_rot~q ),
	.datab(\E_valid_from_R~q ),
	.datac(\E_stall~0_combout ),
	.datad(\E_stall~1_combout ),
	.cin(gnd),
	.combout(\E_stall~2_combout ),
	.cout());
defparam \E_stall~2 .lut_mask = 16'hFFFE;
defparam \E_stall~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.cout());
defparam \D_ctrl_ld_signed~0 .lut_mask = 16'hEFFF;
defparam \D_ctrl_ld_signed~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld~2_combout ),
	.cout());
defparam \D_ctrl_ld~2 .lut_mask = 16'hBFBF;
defparam \D_ctrl_ld~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~3 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(\D_iw[0]~q ),
	.datad(\D_ctrl_ld~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_ld~3_combout ),
	.cout());
defparam \D_ctrl_ld~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_ld~3 .sum_lutc_input = "datac";

dffeas R_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

cycloneive_lcell_comb \av_ld_getting_data~0 (
	.dataa(src0_valid),
	.datab(mem_67_0),
	.datac(src0_valid1),
	.datad(mem_67_01),
	.cin(gnd),
	.combout(\av_ld_getting_data~0_combout ),
	.cout());
defparam \av_ld_getting_data~0 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~1 (
	.dataa(out_valid),
	.datab(mem_67_02),
	.datac(read_latency_shift_reg_02),
	.datad(mem_67_03),
	.cin(gnd),
	.combout(\av_ld_getting_data~1_combout ),
	.cout());
defparam \av_ld_getting_data~1 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~2 (
	.dataa(\av_ld_getting_data~0_combout ),
	.datab(\av_ld_getting_data~1_combout ),
	.datac(src0_valid2),
	.datad(mem_67_04),
	.cin(gnd),
	.combout(\av_ld_getting_data~2_combout ),
	.cout());
defparam \av_ld_getting_data~2 .lut_mask = 16'hEFFF;
defparam \av_ld_getting_data~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~3 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_67_05),
	.datac(read_latency_shift_reg_04),
	.datad(mem_67_06),
	.cin(gnd),
	.combout(\av_ld_getting_data~3_combout ),
	.cout());
defparam \av_ld_getting_data~3 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~4 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_67_07),
	.datac(read_latency_shift_reg_05),
	.datad(mem_67_08),
	.cin(gnd),
	.combout(\av_ld_getting_data~4_combout ),
	.cout());
defparam \av_ld_getting_data~4 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~5 (
	.dataa(\av_ld_getting_data~3_combout ),
	.datab(\av_ld_getting_data~4_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_67),
	.cin(gnd),
	.combout(\av_ld_getting_data~5_combout ),
	.cout());
defparam \av_ld_getting_data~5 .lut_mask = 16'hEFFF;
defparam \av_ld_getting_data~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~7 (
	.dataa(d_read1),
	.datab(WideOr1),
	.datac(\av_ld_getting_data~2_combout ),
	.datad(\av_ld_getting_data~5_combout ),
	.cin(gnd),
	.combout(\av_ld_getting_data~7_combout ),
	.cout());
defparam \av_ld_getting_data~7 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~7 .sum_lutc_input = "datac";

dffeas av_ld_waiting_for_data(
	.clk(clk_clk),
	.d(\av_ld_waiting_for_data_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cycloneive_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(\av_ld_getting_data~7_combout ),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_ld~q ),
	.datad(\av_ld_waiting_for_data~q ),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 16'hFAFC;
defparam \av_ld_waiting_for_data_nxt~0 .sum_lutc_input = "datac";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_aligning_data_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[0]~0 (
	.dataa(\av_ld_align_cycle[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\av_ld_getting_data~7_combout ),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~0_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[0]~0 .lut_mask = 16'hFF55;
defparam \av_ld_align_cycle_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[0] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_mem16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.cout());
defparam \D_ctrl_mem16~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_mem16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem16~1 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.cout());
defparam \D_ctrl_mem16~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[1]~1 (
	.dataa(\av_ld_getting_data~7_combout ),
	.datab(gnd),
	.datac(\av_ld_align_cycle[1]~q ),
	.datad(\av_ld_align_cycle[0]~q ),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~1_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[1]~1 .lut_mask = 16'hAFFA;
defparam \av_ld_align_cycle_nxt[1]~1 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[1] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_align_cycle[0]~q ),
	.datac(\D_ctrl_mem16~1_combout ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 16'hBEFF;
defparam \av_ld_aligning_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem32~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.cout());
defparam \D_ctrl_mem32~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem32~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(\av_ld_aligning_data_nxt~0_combout ),
	.datab(\av_ld_getting_data~7_combout ),
	.datac(\av_ld_aligning_data~q ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 16'hBFFF;
defparam \av_ld_aligning_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~3 (
	.dataa(\E_valid_from_R~q ),
	.datab(\av_ld_waiting_for_data_nxt~0_combout ),
	.datac(\av_ld_aligning_data_nxt~1_combout ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\E_stall~3_combout ),
	.cout());
defparam \E_stall~3 .lut_mask = 16'hFEFF;
defparam \E_stall~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~4 (
	.dataa(\E_stall~2_combout ),
	.datab(\R_ctrl_ld~q ),
	.datac(\E_new_inst~q ),
	.datad(\E_stall~3_combout ),
	.cin(gnd),
	.combout(\E_stall~4_combout ),
	.cout());
defparam \E_stall~4 .lut_mask = 16'hFFFE;
defparam \E_stall~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~3 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\R_valid~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_valid_from_R~3_combout ),
	.cout());
defparam \E_valid_from_R~3 .lut_mask = 16'hFEFE;
defparam \E_valid_from_R~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~2 (
	.dataa(\E_stall~4_combout ),
	.datab(d_write1),
	.datac(av_waitrequest),
	.datad(\E_valid_from_R~3_combout ),
	.cin(gnd),
	.combout(\E_valid_from_R~2_combout ),
	.cout());
defparam \E_valid_from_R~2 .lut_mask = 16'hFFFE;
defparam \E_valid_from_R~2 .sum_lutc_input = "datac";

dffeas E_valid_from_R(
	.clk(clk_clk),
	.d(\E_valid_from_R~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cycloneive_lcell_comb \D_ctrl_jmp_direct~1 (
	.dataa(\D_ctrl_jmp_direct~0_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~1_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_jmp_direct~1 .sum_lutc_input = "datac";

dffeas R_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_direct~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

cycloneive_lcell_comb \R_src1~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_valid_from_R~q ),
	.datad(\R_ctrl_jmp_direct~q ),
	.cin(gnd),
	.combout(\R_src1~10_combout ),
	.cout());
defparam \R_src1~10 .lut_mask = 16'h0FFF;
defparam \R_src1~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[6]~24 (
	.dataa(\D_iw[10]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[6]~24_combout ),
	.cout());
defparam \E_src1[6]~24 .lut_mask = 16'hAACC;
defparam \E_src1[6]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[0]~0 (
	.dataa(F_pc_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\F_pc_plus_one[0]~0_combout ),
	.cout(\F_pc_plus_one[0]~1 ));
defparam \F_pc_plus_one[0]~0 .lut_mask = 16'h55AA;
defparam \F_pc_plus_one[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[1]~2 (
	.dataa(F_pc_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[0]~1 ),
	.combout(\F_pc_plus_one[1]~2_combout ),
	.cout(\F_pc_plus_one[1]~3 ));
defparam \F_pc_plus_one[1]~2 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[2]~4 (
	.dataa(F_pc_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[1]~3 ),
	.combout(\F_pc_plus_one[2]~4_combout ),
	.cout(\F_pc_plus_one[2]~5 ));
defparam \F_pc_plus_one[2]~4 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[3]~6 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[2]~5 ),
	.combout(\F_pc_plus_one[3]~6_combout ),
	.cout(\F_pc_plus_one[3]~7 ));
defparam \F_pc_plus_one[3]~6 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[4]~8 (
	.dataa(F_pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[3]~7 ),
	.combout(\F_pc_plus_one[4]~8_combout ),
	.cout(\F_pc_plus_one[4]~9 ));
defparam \F_pc_plus_one[4]~8 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[4]~8 .sum_lutc_input = "cin";

dffeas R_ctrl_br(
	.clk(clk_clk),
	.d(\R_ctrl_br_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cycloneive_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(\Equal62~9_combout ),
	.datab(\Equal62~12_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.cout());
defparam \D_ctrl_retaddr~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_retaddr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~4 (
	.dataa(\D_ctrl_retaddr~3_combout ),
	.datab(\Equal62~8_combout ),
	.datac(\Equal62~14_combout ),
	.datad(\D_dst_regnum[0]~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~4_combout ),
	.cout());
defparam \D_ctrl_retaddr~4 .lut_mask = 16'hFEFF;
defparam \D_ctrl_retaddr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~5 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_retaddr~4_combout ),
	.datac(\D_ctrl_force_src2_zero~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~5_combout ),
	.cout());
defparam \D_ctrl_retaddr~5 .lut_mask = 16'hF7F7;
defparam \D_ctrl_retaddr~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~9 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hFF7F;
defparam \Equal0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~6 (
	.dataa(\Equal0~12_combout ),
	.datab(\D_ctrl_exception~2_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~6_combout ),
	.cout());
defparam \D_ctrl_retaddr~6 .lut_mask = 16'hFDFE;
defparam \D_ctrl_retaddr~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~7 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~16_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~7_combout ),
	.cout());
defparam \D_ctrl_retaddr~7 .lut_mask = 16'hFFBE;
defparam \D_ctrl_retaddr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~8 (
	.dataa(\Equal0~2_combout ),
	.datab(\D_ctrl_retaddr~5_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~8_combout ),
	.cout());
defparam \D_ctrl_retaddr~8 .lut_mask = 16'hBFFB;
defparam \D_ctrl_retaddr~8 .sum_lutc_input = "datac";

dffeas R_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cycloneive_lcell_comb \R_src1~11 (
	.dataa(\R_valid~q ),
	.datab(\E_valid_from_R~q ),
	.datac(\R_ctrl_br~q ),
	.datad(\R_ctrl_retaddr~q ),
	.cin(gnd),
	.combout(\R_src1~11_combout ),
	.cout());
defparam \R_src1~11 .lut_mask = 16'hFFFE;
defparam \R_src1~11 .sum_lutc_input = "datac";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~24_combout ),
	.asdata(\F_pc_plus_one[4]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cycloneive_lcell_comb D_op_wrctl(
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~3_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_wrctl~combout ),
	.cout());
defparam D_op_wrctl.lut_mask = 16'hFEFF;
defparam D_op_wrctl.sum_lutc_input = "datac";

dffeas R_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cycloneive_lcell_comb \W_ienable_reg_nxt~0 (
	.dataa(\D_iw[7]~q ),
	.datab(\R_ctrl_wrctl_inst~q ),
	.datac(gnd),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~0_combout ),
	.cout());
defparam \W_ienable_reg_nxt~0 .lut_mask = 16'hEEFF;
defparam \W_ienable_reg_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_ienable_reg_nxt~1 (
	.dataa(\E_valid_from_R~q ),
	.datab(\D_iw[6]~q ),
	.datac(\W_ienable_reg_nxt~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~1_combout ),
	.cout());
defparam \W_ienable_reg_nxt~1 .lut_mask = 16'hFEFE;
defparam \W_ienable_reg_nxt~1 .sum_lutc_input = "datac";

dffeas \W_ienable_reg[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~1_combout ),
	.q(\W_ienable_reg[6]~q ),
	.prn(vcc));
defparam \W_ienable_reg[6] .is_wysiwyg = "true";
defparam \W_ienable_reg[6] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[6]~0 (
	.dataa(\W_ienable_reg[6]~q ),
	.datab(dreg_1),
	.datac(gnd),
	.datad(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[6]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[6]~0_combout ),
	.cout());
defparam \W_ipending_reg_nxt[6]~0 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[6]~0 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[6] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[6]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[6]~q ),
	.prn(vcc));
defparam \W_ipending_reg[6] .is_wysiwyg = "true";
defparam \W_ipending_reg[6] .power_up = "low";

cycloneive_lcell_comb \E_src1[5]~25 (
	.dataa(\D_iw[9]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[5]~25_combout ),
	.cout());
defparam \E_src1[5]~25 .lut_mask = 16'hAACC;
defparam \E_src1[5]~25 .sum_lutc_input = "datac";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~25_combout ),
	.asdata(\F_pc_plus_one[3]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

dffeas \W_ienable_reg[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~1_combout ),
	.q(\W_ienable_reg[5]~q ),
	.prn(vcc));
defparam \W_ienable_reg[5] .is_wysiwyg = "true";
defparam \W_ienable_reg[5] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[5]~1 (
	.dataa(\W_ienable_reg[5]~q ),
	.datab(av_readdata_9),
	.datac(av_readdata_8),
	.datad(\the_usb_system_cpu_cpu_nios2_oci|the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[5]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[5]~1_combout ),
	.cout());
defparam \W_ipending_reg_nxt[5]~1 .lut_mask = 16'hFEFF;
defparam \W_ipending_reg_nxt[5]~1 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[5] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[5]~q ),
	.prn(vcc));
defparam \W_ipending_reg[5] .is_wysiwyg = "true";
defparam \W_ipending_reg[5] .power_up = "low";

cycloneive_lcell_comb \R_src1[0]~13 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[0]~13_combout ),
	.cout());
defparam \R_src1[0]~13 .lut_mask = 16'hF7FF;
defparam \R_src1[0]~13 .sum_lutc_input = "datac";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\R_src1[0]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cycloneive_lcell_comb \E_wrctl_estatus~0 (
	.dataa(\D_iw[6]~q ),
	.datab(\R_ctrl_wrctl_inst~q ),
	.datac(\D_iw[8]~q ),
	.datad(\D_iw[7]~q ),
	.cin(gnd),
	.combout(\E_wrctl_estatus~0_combout ),
	.cout());
defparam \E_wrctl_estatus~0 .lut_mask = 16'hEFFF;
defparam \E_wrctl_estatus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~4 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~14_combout ),
	.datac(\Equal62~8_combout ),
	.datad(\D_dst_regnum[0]~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~4_combout ),
	.cout());
defparam \D_ctrl_exception~4 .lut_mask = 16'hFEFF;
defparam \D_ctrl_exception~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~19 (
	.dataa(\D_iw[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~19_combout ),
	.cout());
defparam \D_dst_regnum[0]~19 .lut_mask = 16'hAAFF;
defparam \D_dst_regnum[0]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~5 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~5_combout ),
	.cout());
defparam \D_ctrl_exception~5 .lut_mask = 16'hFBFF;
defparam \D_ctrl_exception~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~6 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_exception~4_combout ),
	.datac(\D_dst_regnum[0]~19_combout ),
	.datad(\D_ctrl_exception~5_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~6_combout ),
	.cout());
defparam \D_ctrl_exception~6 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~0 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~12_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.cout());
defparam \D_ctrl_exception~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_exception~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~1 (
	.dataa(\Equal0~3_combout ),
	.datab(\Equal0~2_combout ),
	.datac(\Equal0~16_combout ),
	.datad(\D_ctrl_exception~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.cout());
defparam \D_ctrl_exception~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~3 (
	.dataa(\D_ctrl_exception~1_combout ),
	.datab(\D_ctrl_exception~2_combout ),
	.datac(\Equal0~12_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~3_combout ),
	.cout());
defparam \D_ctrl_exception~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_exception~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~7 (
	.dataa(\D_ctrl_exception~6_combout ),
	.datab(\D_dst_regnum[0]~21_combout ),
	.datac(\D_dst_regnum[0]~11_combout ),
	.datad(\D_ctrl_exception~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~7_combout ),
	.cout());
defparam \D_ctrl_exception~7 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~7 .sum_lutc_input = "datac";

dffeas R_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_estatus_reg~q ),
	.datac(\E_wrctl_estatus~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 16'hACFF;
defparam \W_estatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~1 (
	.dataa(\W_estatus_reg_inst_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\W_status_reg_pie~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~1 .lut_mask = 16'hFEFE;
defparam \W_estatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_estatus_reg(
	.clk(clk_clk),
	.d(\W_estatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\E_src1[0]~q ),
	.datac(\W_ienable_reg_nxt~0_combout ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 16'hEFFE;
defparam \W_bstatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_break~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\D_iw[16]~q ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.cout());
defparam \D_ctrl_break~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_break~0 .sum_lutc_input = "datac";

dffeas R_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~1 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\W_bstatus_reg_inst_nxt~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~1 .lut_mask = 16'hAACC;
defparam \W_bstatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_bstatus_reg(
	.clk(clk_clk),
	.d(\W_bstatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cycloneive_lcell_comb \E_wrctl_status~0 (
	.dataa(\R_ctrl_wrctl_inst~q ),
	.datab(\D_iw[8]~q ),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~0_combout ),
	.cout());
defparam \E_wrctl_status~0 .lut_mask = 16'hBFFF;
defparam \E_wrctl_status~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_status_reg_pie~q ),
	.datac(gnd),
	.datad(\E_wrctl_status~0_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 16'hAACC;
defparam \W_status_reg_pie_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~0_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\Equal62~10_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_op_eret(
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~10_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_eret~combout ),
	.cout());
defparam D_op_eret.lut_mask = 16'hEFFF;
defparam D_op_eret.sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_sel_nxt.10~1 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\R_ctrl_break~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~1_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~1 .lut_mask = 16'hEEEE;
defparam \F_pc_sel_nxt.10~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(\W_estatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~1_combout ),
	.datac(\D_op_eret~combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 16'hACFF;
defparam \W_status_reg_pie_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cycloneive_lcell_comb \D_iw[5]~0 (
	.dataa(gnd),
	.datab(\W_ipending_reg[6]~q ),
	.datac(\W_ipending_reg[5]~q ),
	.datad(\W_status_reg_pie~q ),
	.cin(gnd),
	.combout(\D_iw[5]~0_combout ),
	.cout());
defparam \D_iw[5]~0 .lut_mask = 16'h3FFF;
defparam \D_iw[5]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_iw[5]~1 (
	.dataa(\D_iw[5]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(gnd),
	.datad(\hbreak_req~0_combout ),
	.cin(gnd),
	.combout(\D_iw[5]~1_combout ),
	.cout());
defparam \D_iw[5]~1 .lut_mask = 16'hEEFF;
defparam \D_iw[5]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[11]~26 (
	.dataa(\F_iw[11]~25_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[11]~26_combout ),
	.cout());
defparam \F_iw[11]~26 .lut_mask = 16'hFEFF;
defparam \F_iw[11]~26 .sum_lutc_input = "datac";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cycloneive_lcell_comb \Equal62~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~0_combout ),
	.cout());
defparam \Equal62~0 .lut_mask = 16'h7FFF;
defparam \Equal62~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hFFBF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~8 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~5_combout ),
	.datad(\D_ctrl_alu_force_xor~14_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~8_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~8 .lut_mask = 16'h27FF;
defparam \D_ctrl_alu_subtract~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~9 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_alu_subtract~8_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~9_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~9 .lut_mask = 16'hEEFF;
defparam \D_ctrl_alu_subtract~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~5 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~5_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~5 .lut_mask = 16'hFF96;
defparam \D_ctrl_alu_subtract~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~10 (
	.dataa(\D_ctrl_alu_subtract~5_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~10_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~10 .lut_mask = 16'hBFBF;
defparam \D_ctrl_alu_subtract~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_alu_sub~0 (
	.dataa(\R_valid~q ),
	.datab(\D_ctrl_alu_subtract~9_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_subtract~10_combout ),
	.cin(gnd),
	.combout(\E_alu_sub~0_combout ),
	.cout());
defparam \E_alu_sub~0 .lut_mask = 16'hFFFE;
defparam \E_alu_sub~0 .sum_lutc_input = "datac";

dffeas E_alu_sub(
	.clk(clk_clk),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cycloneive_lcell_comb \E_src2[12]~15 (
	.dataa(\R_ctrl_src_imm5_shift_rot~q ),
	.datab(\R_ctrl_hi_imm16~q ),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[12]~15_combout ),
	.cout());
defparam \E_src2[12]~15 .lut_mask = 16'hFEFE;
defparam \E_src2[12]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[7]~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[7]~0_combout ),
	.cout());
defparam \R_src2_lo[7]~0 .lut_mask = 16'hACFF;
defparam \R_src2_lo[7]~0 .sum_lutc_input = "datac";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\R_src2_lo[7]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[7]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[7]~23 (
	.dataa(\D_iw[11]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[7]~23_combout ),
	.cout());
defparam \E_src1[7]~23 .lut_mask = 16'hAACC;
defparam \E_src1[7]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[5]~10 (
	.dataa(F_pc_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[4]~9 ),
	.combout(\F_pc_plus_one[5]~10_combout ),
	.cout(\F_pc_plus_one[5]~11 ));
defparam \F_pc_plus_one[5]~10 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[5]~10 .sum_lutc_input = "cin";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\E_src1[7]~23_combout ),
	.asdata(\F_pc_plus_one[5]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[6]~1 (
	.dataa(\D_iw[12]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[6]~1_combout ),
	.cout());
defparam \R_src2_lo[6]~1 .lut_mask = 16'hACFF;
defparam \R_src2_lo[6]~1 .sum_lutc_input = "datac";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\R_src2_lo[6]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[6]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[5]~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[5]~2_combout ),
	.cout());
defparam \R_src2_lo[5]~2 .lut_mask = 16'hACFF;
defparam \R_src2_lo[5]~2 .sum_lutc_input = "datac";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\R_src2_lo[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[5]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_src2[4]~q ),
	.datad(\E_alu_sub~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[4]~26 (
	.dataa(\D_iw[8]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[4]~26_combout ),
	.cout());
defparam \E_src1[4]~26 .lut_mask = 16'hAACC;
defparam \E_src1[4]~26 .sum_lutc_input = "datac";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\E_src1[4]~26_combout ),
	.asdata(\F_pc_plus_one[2]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[3]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[3]~8 (
	.dataa(\D_iw[7]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[3]~8_combout ),
	.cout());
defparam \E_src1[3]~8 .lut_mask = 16'hAACC;
defparam \E_src1[3]~8 .sum_lutc_input = "datac";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\E_src1[3]~8_combout ),
	.asdata(\F_pc_plus_one[1]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cycloneive_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[2]~q ),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[2]~7 (
	.dataa(\D_iw[6]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[2]~7_combout ),
	.cout());
defparam \E_src1[2]~7 .lut_mask = 16'hAACC;
defparam \E_src1[2]~7 .sum_lutc_input = "datac";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\E_src1[2]~7_combout ),
	.asdata(\F_pc_plus_one[0]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[1]~q ),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[1]~12 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[1]~12_combout ),
	.cout());
defparam \R_src1[1]~12 .lut_mask = 16'hF7FF;
defparam \R_src1[1]~12 .sum_lutc_input = "datac";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\R_src1[1]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

cycloneive_lcell_comb \Add1~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[0]~q ),
	.cin(gnd),
	.combout(\Add1~7_combout ),
	.cout());
defparam \Add1~7 .lut_mask = 16'h0FF0;
defparam \Add1~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~9 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add1~9_cout ));
defparam \Add1~9 .lut_mask = 16'h00AA;
defparam \Add1~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~10 (
	.dataa(\Add1~7_combout ),
	.datab(\E_src1[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9_cout ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
defparam \Add1~10 .lut_mask = 16'h967F;
defparam \Add1~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~12 (
	.dataa(\Add1~6_combout ),
	.datab(\E_src1[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
defparam \Add1~12 .lut_mask = 16'h96EF;
defparam \Add1~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~14 (
	.dataa(\Add1~5_combout ),
	.datab(\E_src1[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
defparam \Add1~14 .lut_mask = 16'h967F;
defparam \Add1~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~16 (
	.dataa(\Add1~4_combout ),
	.datab(\E_src1[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
defparam \Add1~16 .lut_mask = 16'h96EF;
defparam \Add1~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~18 (
	.dataa(\Add1~3_combout ),
	.datab(\E_src1[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
defparam \Add1~18 .lut_mask = 16'h967F;
defparam \Add1~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~20 (
	.dataa(\Add1~2_combout ),
	.datab(\E_src1[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
defparam \Add1~20 .lut_mask = 16'h96EF;
defparam \Add1~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~22 (
	.dataa(\Add1~1_combout ),
	.datab(\E_src1[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
defparam \Add1~22 .lut_mask = 16'h967F;
defparam \Add1~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~24 (
	.dataa(\Add1~0_combout ),
	.datab(\E_src1[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
defparam \Add1~24 .lut_mask = 16'h96EF;
defparam \Add1~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.cout());
defparam \D_logic_op_raw[1]~0 .lut_mask = 16'hEFFF;
defparam \D_logic_op_raw[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~10 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(\D_ctrl_alu_force_xor~14_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~10_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~10 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~11 (
	.dataa(\Equal0~5_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~11_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~11 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~13 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~13_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~13 .lut_mask = 16'hFFD8;
defparam \D_ctrl_alu_force_xor~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~12 (
	.dataa(\D_ctrl_alu_force_xor~10_combout ),
	.datab(\D_ctrl_alu_force_xor~11_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_force_xor~13_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~12_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~12 .lut_mask = 16'hFFFE;
defparam \D_ctrl_alu_force_xor~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_logic_op[1]~0 (
	.dataa(\D_logic_op_raw[1]~0_combout ),
	.datab(\D_ctrl_alu_force_xor~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.cout());
defparam \D_logic_op[1]~0 .lut_mask = 16'hEEEE;
defparam \D_logic_op[1]~0 .sum_lutc_input = "datac";

dffeas \R_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op[0]~1 (
	.dataa(\D_ctrl_alu_force_xor~12_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\Equal0~7_combout ),
	.cin(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.cout());
defparam \D_logic_op[0]~1 .lut_mask = 16'hFAFC;
defparam \D_logic_op[0]~1 .sum_lutc_input = "datac";

dffeas \R_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[7]~0 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[7]~q ),
	.datac(\E_src1[7]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[7]~0_combout ),
	.cout());
defparam \E_logic_result[7]~0 .lut_mask = 16'h6996;
defparam \E_logic_result[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~8 (
	.dataa(\D_iw[13]~q ),
	.datab(gnd),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'hAFFF;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~10 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
defparam \Equal0~10 .lut_mask = 16'hFFF7;
defparam \Equal0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_logic~0 (
	.dataa(gnd),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~9_combout ),
	.datad(\Equal0~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.cout());
defparam \D_ctrl_logic~0 .lut_mask = 16'h3FFF;
defparam \D_ctrl_logic~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_ctrl_logic(
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\Equal0~8_combout ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~combout ),
	.cout());
defparam D_ctrl_logic.lut_mask = 16'hFEFF;
defparam D_ctrl_logic.sum_lutc_input = "datac";

dffeas R_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cycloneive_lcell_comb \W_alu_result[7]~23 (
	.dataa(\Add1~24_combout ),
	.datab(\E_logic_result[7]~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[7]~23_combout ),
	.cout());
defparam \W_alu_result[7]~23 .lut_mask = 16'hAACC;
defparam \W_alu_result[7]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_shift_rot_right~0_combout ),
	.datad(\D_iw[13]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~1 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[6]~14 (
	.dataa(\E_shift_rot_result[7]~q ),
	.datab(\E_shift_rot_result[5]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[6]~14_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[6]~14 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[6]~14 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[6]~14_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[5]~24 (
	.dataa(\E_shift_rot_result[6]~q ),
	.datab(\E_shift_rot_result[4]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[5]~24_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[5]~24 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[5]~24 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[5]~24_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[4]~23 (
	.dataa(\E_shift_rot_result[5]~q ),
	.datab(\E_shift_rot_result[3]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[4]~23_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[4]~23 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[4]~23 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[4]~23_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[3]~26 (
	.dataa(\E_shift_rot_result[4]~q ),
	.datab(\E_shift_rot_result[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[3]~26_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[3]~26 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[3]~26 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[3]~26_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[2]~25 (
	.dataa(\E_shift_rot_result[3]~q ),
	.datab(\E_shift_rot_result[1]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[2]~25_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[2]~25 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[2]~25 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[2]~25_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[1]~28 (
	.dataa(\E_shift_rot_result[2]~q ),
	.datab(\E_shift_rot_result[0]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[1]~28_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[1]~28 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[1]~28 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[1]~28_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[0]~29 (
	.dataa(\E_shift_rot_result[1]~q ),
	.datab(\E_shift_rot_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[0]~29_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[0]~29 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[0]~29 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[0]~29_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cycloneive_lcell_comb \R_ctrl_rot_right_nxt~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~7_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\R_ctrl_rot_right_nxt~0_combout ),
	.cout());
defparam \R_ctrl_rot_right_nxt~0 .lut_mask = 16'hFEFF;
defparam \R_ctrl_rot_right_nxt~0 .sum_lutc_input = "datac";

dffeas R_ctrl_rot_right(
	.clk(clk_clk),
	.d(\R_ctrl_rot_right_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cycloneive_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~4_combout ),
	.datad(\Equal62~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.cout());
defparam \D_ctrl_shift_logical~1 .lut_mask = 16'hFFB8;
defparam \D_ctrl_shift_logical~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[15]~q ),
	.datac(\D_ctrl_shift_logical~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~2_combout ),
	.cout());
defparam \D_ctrl_shift_logical~2 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_logical~2 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(\E_shift_rot_result[0]~q ),
	.datab(\E_shift_rot_result[31]~q ),
	.datac(\R_ctrl_rot_right~q ),
	.datad(\R_ctrl_shift_logical~q ),
	.cin(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.cout());
defparam \E_shift_rot_fill_bit~0 .lut_mask = 16'hACFF;
defparam \E_shift_rot_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_result_nxt[31]~31 (
	.dataa(\E_shift_rot_fill_bit~0_combout ),
	.datab(\E_shift_rot_result[30]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[31]~31_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[31]~31 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[31]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[31]~14 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[31]~14_combout ),
	.cout());
defparam \R_src1[31]~14 .lut_mask = 16'hF7FF;
defparam \R_src1[31]~14 .sum_lutc_input = "datac";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\R_src1[31]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[31]~31_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[30]~30 (
	.dataa(\E_shift_rot_result[31]~q ),
	.datab(\E_shift_rot_result[29]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[30]~30_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[30]~30 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[30]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[30]~16 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[30]~16_combout ),
	.cout());
defparam \R_src1[30]~16 .lut_mask = 16'hF7FF;
defparam \R_src1[30]~16 .sum_lutc_input = "datac";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\R_src1[30]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[30]~30_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[29]~27 (
	.dataa(\E_shift_rot_result[30]~q ),
	.datab(\E_shift_rot_result[28]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[29]~27_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[29]~27 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[29]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[29]~15 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[29]~15_combout ),
	.cout());
defparam \R_src1[29]~15 .lut_mask = 16'hF7FF;
defparam \R_src1[29]~15 .sum_lutc_input = "datac";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\R_src1[29]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[29]~27_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[28]~19 (
	.dataa(\E_shift_rot_result[29]~q ),
	.datab(\E_shift_rot_result[27]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[28]~19_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[28]~19 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[28]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[28]~0 (
	.dataa(F_pc_26),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[28]~0_combout ),
	.cout());
defparam \E_src1[28]~0 .lut_mask = 16'hAACC;
defparam \E_src1[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[6]~12 (
	.dataa(F_pc_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[5]~11 ),
	.combout(\F_pc_plus_one[6]~12_combout ),
	.cout(\F_pc_plus_one[6]~13 ));
defparam \F_pc_plus_one[6]~12 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[7]~14 (
	.dataa(F_pc_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[6]~13 ),
	.combout(\F_pc_plus_one[7]~14_combout ),
	.cout(\F_pc_plus_one[7]~15 ));
defparam \F_pc_plus_one[7]~14 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[8]~16 (
	.dataa(F_pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[7]~15 ),
	.combout(\F_pc_plus_one[8]~16_combout ),
	.cout(\F_pc_plus_one[8]~17 ));
defparam \F_pc_plus_one[8]~16 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[9]~18 (
	.dataa(F_pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[8]~17 ),
	.combout(\F_pc_plus_one[9]~18_combout ),
	.cout(\F_pc_plus_one[9]~19 ));
defparam \F_pc_plus_one[9]~18 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[9]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[10]~20 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[9]~19 ),
	.combout(\F_pc_plus_one[10]~20_combout ),
	.cout(\F_pc_plus_one[10]~21 ));
defparam \F_pc_plus_one[10]~20 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[10]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[11]~22 (
	.dataa(F_pc_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[10]~21 ),
	.combout(\F_pc_plus_one[11]~22_combout ),
	.cout(\F_pc_plus_one[11]~23 ));
defparam \F_pc_plus_one[11]~22 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[11]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[12]~24 (
	.dataa(F_pc_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[11]~23 ),
	.combout(\F_pc_plus_one[12]~24_combout ),
	.cout(\F_pc_plus_one[12]~25 ));
defparam \F_pc_plus_one[12]~24 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[12]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[13]~26 (
	.dataa(F_pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[12]~25 ),
	.combout(\F_pc_plus_one[13]~26_combout ),
	.cout(\F_pc_plus_one[13]~27 ));
defparam \F_pc_plus_one[13]~26 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[13]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[14]~28 (
	.dataa(F_pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[13]~27 ),
	.combout(\F_pc_plus_one[14]~28_combout ),
	.cout(\F_pc_plus_one[14]~29 ));
defparam \F_pc_plus_one[14]~28 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[14]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[15]~30 (
	.dataa(F_pc_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[14]~29 ),
	.combout(\F_pc_plus_one[15]~30_combout ),
	.cout(\F_pc_plus_one[15]~31 ));
defparam \F_pc_plus_one[15]~30 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[15]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[16]~32 (
	.dataa(F_pc_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[15]~31 ),
	.combout(\F_pc_plus_one[16]~32_combout ),
	.cout(\F_pc_plus_one[16]~33 ));
defparam \F_pc_plus_one[16]~32 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[16]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[17]~34 (
	.dataa(F_pc_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[16]~33 ),
	.combout(\F_pc_plus_one[17]~34_combout ),
	.cout(\F_pc_plus_one[17]~35 ));
defparam \F_pc_plus_one[17]~34 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[17]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[18]~36 (
	.dataa(F_pc_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[17]~35 ),
	.combout(\F_pc_plus_one[18]~36_combout ),
	.cout(\F_pc_plus_one[18]~37 ));
defparam \F_pc_plus_one[18]~36 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[18]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[19]~38 (
	.dataa(F_pc_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[18]~37 ),
	.combout(\F_pc_plus_one[19]~38_combout ),
	.cout(\F_pc_plus_one[19]~39 ));
defparam \F_pc_plus_one[19]~38 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[19]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[20]~40 (
	.dataa(F_pc_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[19]~39 ),
	.combout(\F_pc_plus_one[20]~40_combout ),
	.cout(\F_pc_plus_one[20]~41 ));
defparam \F_pc_plus_one[20]~40 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[20]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[21]~42 (
	.dataa(F_pc_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[20]~41 ),
	.combout(\F_pc_plus_one[21]~42_combout ),
	.cout(\F_pc_plus_one[21]~43 ));
defparam \F_pc_plus_one[21]~42 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[21]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[22]~44 (
	.dataa(F_pc_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[21]~43 ),
	.combout(\F_pc_plus_one[22]~44_combout ),
	.cout(\F_pc_plus_one[22]~45 ));
defparam \F_pc_plus_one[22]~44 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[22]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[23]~46 (
	.dataa(F_pc_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[22]~45 ),
	.combout(\F_pc_plus_one[23]~46_combout ),
	.cout(\F_pc_plus_one[23]~47 ));
defparam \F_pc_plus_one[23]~46 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[23]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[24]~48 (
	.dataa(F_pc_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[23]~47 ),
	.combout(\F_pc_plus_one[24]~48_combout ),
	.cout(\F_pc_plus_one[24]~49 ));
defparam \F_pc_plus_one[24]~48 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[24]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[25]~50 (
	.dataa(F_pc_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[24]~49 ),
	.combout(\F_pc_plus_one[25]~50_combout ),
	.cout(\F_pc_plus_one[25]~51 ));
defparam \F_pc_plus_one[25]~50 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[25]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[26]~52 (
	.dataa(F_pc_26),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\F_pc_plus_one[25]~51 ),
	.combout(\F_pc_plus_one[26]~52_combout ),
	.cout());
defparam \F_pc_plus_one[26]~52 .lut_mask = 16'h5A5A;
defparam \F_pc_plus_one[26]~52 .sum_lutc_input = "cin";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\E_src1[28]~0_combout ),
	.asdata(\F_pc_plus_one[26]~52_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

dffeas \E_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[28]~19_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[27]~20 (
	.dataa(\E_shift_rot_result[28]~q ),
	.datab(\E_shift_rot_result[26]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[27]~20_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[27]~20 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[27]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~58 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\F_iw[31]~58_combout ),
	.cout());
defparam \F_iw[31]~58 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~59 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[31]~58_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_31),
	.cin(gnd),
	.combout(\F_iw[31]~59_combout ),
	.cout());
defparam \F_iw[31]~59 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~59 .sum_lutc_input = "datac";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~59_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cycloneive_lcell_comb \E_src1[27]~1 (
	.dataa(\D_iw[31]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[27]~1_combout ),
	.cout());
defparam \E_src1[27]~1 .lut_mask = 16'hAACC;
defparam \E_src1[27]~1 .sum_lutc_input = "datac";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\E_src1[27]~1_combout ),
	.asdata(\F_pc_plus_one[25]~50_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

dffeas \E_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[27]~20_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[26]~21 (
	.dataa(\E_shift_rot_result[27]~q ),
	.datab(\E_shift_rot_result[25]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[26]~21_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[26]~21 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[26]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~60 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_30),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\F_iw[30]~60_combout ),
	.cout());
defparam \F_iw[30]~60 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~61 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[30]~60_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[30]~61_combout ),
	.cout());
defparam \F_iw[30]~61 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~61 .sum_lutc_input = "datac";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~61_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

cycloneive_lcell_comb \E_src1[26]~2 (
	.dataa(\D_iw[30]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[26]~2_combout ),
	.cout());
defparam \E_src1[26]~2 .lut_mask = 16'hAACC;
defparam \E_src1[26]~2 .sum_lutc_input = "datac";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\E_src1[26]~2_combout ),
	.asdata(\F_pc_plus_one[24]~48_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

dffeas \E_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[26]~21_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[25]~22 (
	.dataa(\E_shift_rot_result[26]~q ),
	.datab(\E_shift_rot_result[24]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[25]~22_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[25]~22 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[25]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~62 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_29),
	.cin(gnd),
	.combout(\F_iw[29]~62_combout ),
	.cout());
defparam \F_iw[29]~62 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~63 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[29]~62_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_29),
	.cin(gnd),
	.combout(\F_iw[29]~63_combout ),
	.cout());
defparam \F_iw[29]~63 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~63 .sum_lutc_input = "datac";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~63_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

cycloneive_lcell_comb \E_src1[25]~3 (
	.dataa(\D_iw[29]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[25]~3_combout ),
	.cout());
defparam \E_src1[25]~3 .lut_mask = 16'hAACC;
defparam \E_src1[25]~3 .sum_lutc_input = "datac";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\E_src1[25]~3_combout ),
	.asdata(\F_pc_plus_one[23]~46_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

dffeas \E_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[25]~22_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[24]~15 (
	.dataa(\E_shift_rot_result[25]~q ),
	.datab(\E_shift_rot_result[23]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[24]~15_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[24]~15 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[24]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~56 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_28),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\F_iw[28]~56_combout ),
	.cout());
defparam \F_iw[28]~56 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~57 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[28]~56_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[28]~57_combout ),
	.cout());
defparam \F_iw[28]~57 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~57 .sum_lutc_input = "datac";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~57_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

cycloneive_lcell_comb \E_src1[24]~4 (
	.dataa(\D_iw[28]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[24]~4_combout ),
	.cout());
defparam \E_src1[24]~4 .lut_mask = 16'hAACC;
defparam \E_src1[24]~4 .sum_lutc_input = "datac";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\E_src1[24]~4_combout ),
	.asdata(\F_pc_plus_one[22]~44_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

dffeas \E_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[24]~15_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[23]~11 (
	.dataa(\E_shift_rot_result[24]~q ),
	.datab(\E_shift_rot_result[22]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[23]~11_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[23]~11 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[23]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~54 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_27),
	.cin(gnd),
	.combout(\F_iw[27]~54_combout ),
	.cout());
defparam \F_iw[27]~54 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~55 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[27]~54_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_27),
	.cin(gnd),
	.combout(\F_iw[27]~55_combout ),
	.cout());
defparam \F_iw[27]~55 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~55 .sum_lutc_input = "datac";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~55_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cycloneive_lcell_comb \E_src1[23]~5 (
	.dataa(\D_iw[27]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[23]~5_combout ),
	.cout());
defparam \E_src1[23]~5 .lut_mask = 16'hAACC;
defparam \E_src1[23]~5 .sum_lutc_input = "datac";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\E_src1[23]~5_combout ),
	.asdata(\F_pc_plus_one[21]~42_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

dffeas \E_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[23]~11_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[22]~12 (
	.dataa(\E_shift_rot_result[23]~q ),
	.datab(\E_shift_rot_result[21]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[22]~12_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[22]~12 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[22]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~23 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_26),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\F_iw[26]~23_combout ),
	.cout());
defparam \F_iw[26]~23 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~24 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[26]~23_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[26]~24_combout ),
	.cout());
defparam \F_iw[26]~24 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~24 .sum_lutc_input = "datac";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cycloneive_lcell_comb \E_src1[22]~6 (
	.dataa(\D_iw[26]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[22]~6_combout ),
	.cout());
defparam \E_src1[22]~6 .lut_mask = 16'hAACC;
defparam \E_src1[22]~6 .sum_lutc_input = "datac";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\E_src1[22]~6_combout ),
	.asdata(\F_pc_plus_one[20]~40_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

dffeas \E_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[22]~12_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[21]~16 (
	.dataa(\E_shift_rot_result[22]~q ),
	.datab(\E_shift_rot_result[20]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[21]~16_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[21]~16 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[21]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~21 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\F_iw[25]~21_combout ),
	.cout());
defparam \F_iw[25]~21 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~22 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[25]~21_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_25),
	.cin(gnd),
	.combout(\F_iw[25]~22_combout ),
	.cout());
defparam \F_iw[25]~22 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~22 .sum_lutc_input = "datac";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cycloneive_lcell_comb \E_src1[21]~9 (
	.dataa(\D_iw[25]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[21]~9_combout ),
	.cout());
defparam \E_src1[21]~9 .lut_mask = 16'hAACC;
defparam \E_src1[21]~9 .sum_lutc_input = "datac";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\E_src1[21]~9_combout ),
	.asdata(\F_pc_plus_one[19]~38_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

dffeas \E_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[21]~16_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[20]~17 (
	.dataa(\E_shift_rot_result[21]~q ),
	.datab(\E_shift_rot_result[19]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[20]~17_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[20]~17 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[20]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~19 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_24),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\F_iw[24]~19_combout ),
	.cout());
defparam \F_iw[24]~19 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~20 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[24]~19_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[24]~20_combout ),
	.cout());
defparam \F_iw[24]~20 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~20 .sum_lutc_input = "datac";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cycloneive_lcell_comb \E_src1[20]~10 (
	.dataa(\D_iw[24]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[20]~10_combout ),
	.cout());
defparam \E_src1[20]~10 .lut_mask = 16'hAACC;
defparam \E_src1[20]~10 .sum_lutc_input = "datac";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\E_src1[20]~10_combout ),
	.asdata(\F_pc_plus_one[18]~36_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

dffeas \E_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[20]~17_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[19]~18 (
	.dataa(\E_shift_rot_result[20]~q ),
	.datab(\E_shift_rot_result[18]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[19]~18_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[19]~18 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[19]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~17 (
	.dataa(read_latency_shift_reg_03),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\F_iw[23]~17_combout ),
	.cout());
defparam \F_iw[23]~17 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~18 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[23]~17_combout ),
	.datac(out_valid2),
	.datad(out_data_buffer_23),
	.cin(gnd),
	.combout(\F_iw[23]~18_combout ),
	.cout());
defparam \F_iw[23]~18 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~18 .sum_lutc_input = "datac";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cycloneive_lcell_comb \E_src1[19]~11 (
	.dataa(\D_iw[23]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[19]~11_combout ),
	.cout());
defparam \E_src1[19]~11 .lut_mask = 16'hAACC;
defparam \E_src1[19]~11 .sum_lutc_input = "datac";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\E_src1[19]~11_combout ),
	.asdata(\F_pc_plus_one[17]~34_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

dffeas \E_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[19]~18_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[18]~3 (
	.dataa(\E_shift_rot_result[19]~q ),
	.datab(\E_shift_rot_result[17]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[18]~3_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[18]~3 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[18]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~15 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_22),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\F_iw[22]~15_combout ),
	.cout());
defparam \F_iw[22]~15 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~16 (
	.dataa(\D_iw[5]~1_combout ),
	.datab(\F_iw[22]~15_combout ),
	.datac(src_payload1),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[22]~16_combout ),
	.cout());
defparam \F_iw[22]~16 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~16 .sum_lutc_input = "datac";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cycloneive_lcell_comb \E_src1[18]~12 (
	.dataa(\D_iw[22]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[18]~12_combout ),
	.cout());
defparam \E_src1[18]~12 .lut_mask = 16'hAACC;
defparam \E_src1[18]~12 .sum_lutc_input = "datac";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\E_src1[18]~12_combout ),
	.asdata(\F_pc_plus_one[16]~32_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

dffeas \E_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[18]~3_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[17]~4 (
	.dataa(\E_shift_rot_result[18]~q ),
	.datab(\E_shift_rot_result[16]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[17]~4_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[17]~4 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[17]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[21]~53 (
	.dataa(src_payload5),
	.datab(src1_valid),
	.datac(av_readdata_pre_21),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[21]~53_combout ),
	.cout());
defparam \F_iw[21]~53 .lut_mask = 16'hFEFF;
defparam \F_iw[21]~53 .sum_lutc_input = "datac";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~53_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cycloneive_lcell_comb \E_src1[17]~13 (
	.dataa(\D_iw[21]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[17]~13_combout ),
	.cout());
defparam \E_src1[17]~13 .lut_mask = 16'hAACC;
defparam \E_src1[17]~13 .sum_lutc_input = "datac";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\E_src1[17]~13_combout ),
	.asdata(\F_pc_plus_one[15]~30_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

dffeas \E_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[17]~4_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[16]~5 (
	.dataa(\E_shift_rot_result[17]~q ),
	.datab(\E_shift_rot_result[15]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[16]~5_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[16]~5 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[16]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~47 (
	.dataa(src_payload4),
	.datab(src1_valid),
	.datac(av_readdata_pre_20),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[20]~47_combout ),
	.cout());
defparam \F_iw[20]~47 .lut_mask = 16'hFEFF;
defparam \F_iw[20]~47 .sum_lutc_input = "datac";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cycloneive_lcell_comb \E_src1[16]~14 (
	.dataa(\D_iw[20]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[16]~14_combout ),
	.cout());
defparam \E_src1[16]~14 .lut_mask = 16'hAACC;
defparam \E_src1[16]~14 .sum_lutc_input = "datac";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\E_src1[16]~14_combout ),
	.asdata(\F_pc_plus_one[14]~28_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \E_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[16]~5_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[15]~6 (
	.dataa(\E_shift_rot_result[16]~q ),
	.datab(\E_shift_rot_result[14]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[15]~6_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[15]~6 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[15]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~49 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_19),
	.datad(av_readdata_pre_19),
	.cin(gnd),
	.combout(\F_iw[19]~49_combout ),
	.cout());
defparam \F_iw[19]~49 .lut_mask = 16'hFFFE;
defparam \F_iw[19]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~50 (
	.dataa(\F_iw[19]~49_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(\D_iw[5]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[19]~50_combout ),
	.cout());
defparam \F_iw[19]~50 .lut_mask = 16'hFEFF;
defparam \F_iw[19]~50 .sum_lutc_input = "datac";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cycloneive_lcell_comb \E_src1[15]~15 (
	.dataa(\D_iw[19]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[15]~15_combout ),
	.cout());
defparam \E_src1[15]~15 .lut_mask = 16'hAACC;
defparam \E_src1[15]~15 .sum_lutc_input = "datac";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\E_src1[15]~15_combout ),
	.asdata(\F_pc_plus_one[13]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

dffeas \E_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[15]~6_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[14]~1 (
	.dataa(\E_shift_rot_result[15]~q ),
	.datab(\E_shift_rot_result[13]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[14]~1_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[14]~1 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[14]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~48 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_18),
	.datad(av_readdata_pre_18),
	.cin(gnd),
	.combout(\F_iw[18]~48_combout ),
	.cout());
defparam \F_iw[18]~48 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~65 (
	.dataa(\D_iw[5]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[18]~48_combout ),
	.cin(gnd),
	.combout(\F_iw[18]~65_combout ),
	.cout());
defparam \F_iw[18]~65 .lut_mask = 16'hFFFB;
defparam \F_iw[18]~65 .sum_lutc_input = "datac";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~65_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cycloneive_lcell_comb \E_src1[14]~16 (
	.dataa(\D_iw[18]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[14]~16_combout ),
	.cout());
defparam \E_src1[14]~16 .lut_mask = 16'hAACC;
defparam \E_src1[14]~16 .sum_lutc_input = "datac";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\E_src1[14]~16_combout ),
	.asdata(\F_pc_plus_one[12]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

dffeas \E_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[14]~1_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[13]~2 (
	.dataa(\E_shift_rot_result[14]~q ),
	.datab(\E_shift_rot_result[12]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[13]~2_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[13]~2 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[13]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~51 (
	.dataa(src1_valid),
	.datab(out_valid2),
	.datac(out_data_buffer_17),
	.datad(av_readdata_pre_17),
	.cin(gnd),
	.combout(\F_iw[17]~51_combout ),
	.cout());
defparam \F_iw[17]~51 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~52 (
	.dataa(\F_iw[17]~51_combout ),
	.datab(src_payload1),
	.datac(av_readdata_pre_30),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[17]~52_combout ),
	.cout());
defparam \F_iw[17]~52 .lut_mask = 16'hFEFE;
defparam \F_iw[17]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~66 (
	.dataa(\D_iw[5]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[17]~52_combout ),
	.cin(gnd),
	.combout(\F_iw[17]~66_combout ),
	.cout());
defparam \F_iw[17]~66 .lut_mask = 16'hFFDF;
defparam \F_iw[17]~66 .sum_lutc_input = "datac";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~66_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cycloneive_lcell_comb \E_src1[13]~17 (
	.dataa(\D_iw[17]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[13]~17_combout ),
	.cout());
defparam \E_src1[13]~17 .lut_mask = 16'hAACC;
defparam \E_src1[13]~17 .sum_lutc_input = "datac";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\E_src1[13]~17_combout ),
	.asdata(\F_pc_plus_one[11]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

dffeas \E_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[13]~2_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[12]~7 (
	.dataa(\E_shift_rot_result[13]~q ),
	.datab(\E_shift_rot_result[11]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[12]~7_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[12]~7 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[12]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[12]~18 (
	.dataa(\D_iw[16]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[12]~18_combout ),
	.cout());
defparam \E_src1[12]~18 .lut_mask = 16'hAACC;
defparam \E_src1[12]~18 .sum_lutc_input = "datac";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\E_src1[12]~18_combout ),
	.asdata(\F_pc_plus_one[10]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

dffeas \E_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[12]~7_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[11]~8 (
	.dataa(\E_shift_rot_result[12]~q ),
	.datab(\E_shift_rot_result[10]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[11]~8_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[11]~8 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[11]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[11]~19 (
	.dataa(\D_iw[15]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[11]~19_combout ),
	.cout());
defparam \E_src1[11]~19 .lut_mask = 16'hAACC;
defparam \E_src1[11]~19 .sum_lutc_input = "datac";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\E_src1[11]~19_combout ),
	.asdata(\F_pc_plus_one[9]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

dffeas \E_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[11]~8_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[10]~9 (
	.dataa(\E_shift_rot_result[11]~q ),
	.datab(\E_shift_rot_result[9]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[10]~9_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[10]~9 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[10]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[10]~20 (
	.dataa(\D_iw[14]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[10]~20_combout ),
	.cout());
defparam \E_src1[10]~20 .lut_mask = 16'hAACC;
defparam \E_src1[10]~20 .sum_lutc_input = "datac";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\E_src1[10]~20_combout ),
	.asdata(\F_pc_plus_one[8]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

dffeas \E_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[10]~9_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[9]~10 (
	.dataa(\E_shift_rot_result[10]~q ),
	.datab(\E_shift_rot_result[8]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[9]~10_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[9]~10 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[9]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[9]~21 (
	.dataa(\D_iw[13]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[9]~21_combout ),
	.cout());
defparam \E_src1[9]~21 .lut_mask = 16'hAACC;
defparam \E_src1[9]~21 .sum_lutc_input = "datac";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\E_src1[9]~21_combout ),
	.asdata(\F_pc_plus_one[7]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

dffeas \E_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[9]~10_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[8]~13 (
	.dataa(\E_shift_rot_result[9]~q ),
	.datab(\E_shift_rot_result[7]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[8]~13_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[8]~13 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[8]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[8]~22 (
	.dataa(\D_iw[12]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[8]~22_combout ),
	.cout());
defparam \E_src1[8]~22 .lut_mask = 16'hAACC;
defparam \E_src1[8]~22 .sum_lutc_input = "datac";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\E_src1[8]~22_combout ),
	.asdata(\F_pc_plus_one[6]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

dffeas \E_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[8]~13_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[7]~0 (
	.dataa(\E_shift_rot_result[8]~q ),
	.datab(\E_shift_rot_result[6]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[7]~0_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[7]~0 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[7]~0 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[7]~0_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cycloneive_lcell_comb D_op_rdctl(
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_rdctl~combout ),
	.cout());
defparam D_op_rdctl.lut_mask = 16'hEFFF;
defparam D_op_rdctl.sum_lutc_input = "datac";

dffeas R_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hF7FF;
defparam \Equal0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~2 (
	.dataa(\Equal0~6_combout ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~3_combout ),
	.datad(\D_ctrl_jmp_direct~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~2_combout ),
	.cout());
defparam \D_ctrl_br_cmp~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_br_cmp~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~5 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~5_combout ),
	.cout());
defparam \D_ctrl_br_cmp~5 .lut_mask = 16'hF7B3;
defparam \D_ctrl_br_cmp~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~3 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\D_ctrl_br_cmp~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~3_combout ),
	.cout());
defparam \D_ctrl_br_cmp~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_br_cmp~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~4 (
	.dataa(\D_ctrl_br_cmp~2_combout ),
	.datab(\D_ctrl_br_cmp~3_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~4_combout ),
	.cout());
defparam \D_ctrl_br_cmp~4 .lut_mask = 16'hFFFE;
defparam \D_ctrl_br_cmp~4 .sum_lutc_input = "datac";

dffeas R_ctrl_br_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_br_cmp~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cycloneive_lcell_comb \E_alu_result~0 (
	.dataa(\R_ctrl_rd_ctl_reg~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_alu_result~0_combout ),
	.cout());
defparam \E_alu_result~0 .lut_mask = 16'hEEEE;
defparam \E_alu_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[14]~9 (
	.dataa(\D_iw[20]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[14]~9_combout ),
	.cout());
defparam \R_src2_lo[14]~9 .lut_mask = 16'hACFF;
defparam \R_src2_lo[14]~9 .sum_lutc_input = "datac";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\R_src2_lo[14]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cycloneive_lcell_comb \Add1~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[14]~q ),
	.cin(gnd),
	.combout(\Add1~26_combout ),
	.cout());
defparam \Add1~26 .lut_mask = 16'h0FF0;
defparam \Add1~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[13]~10 (
	.dataa(\D_iw[19]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[13]~10_combout ),
	.cout());
defparam \R_src2_lo[13]~10 .lut_mask = 16'hACFF;
defparam \R_src2_lo[13]~10 .sum_lutc_input = "datac";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\R_src2_lo[13]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cycloneive_lcell_comb \Add1~27 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[13]~q ),
	.cin(gnd),
	.combout(\Add1~27_combout ),
	.cout());
defparam \Add1~27 .lut_mask = 16'h0FF0;
defparam \Add1~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[12]~11 (
	.dataa(\D_iw[18]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[12]~11_combout ),
	.cout());
defparam \R_src2_lo[12]~11 .lut_mask = 16'hACFF;
defparam \R_src2_lo[12]~11 .sum_lutc_input = "datac";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\R_src2_lo[12]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cycloneive_lcell_comb \Add1~28 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[12]~q ),
	.cin(gnd),
	.combout(\Add1~28_combout ),
	.cout());
defparam \Add1~28 .lut_mask = 16'h0FF0;
defparam \Add1~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[11]~12 (
	.dataa(\D_iw[17]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[11]~12_combout ),
	.cout());
defparam \R_src2_lo[11]~12 .lut_mask = 16'hACFF;
defparam \R_src2_lo[11]~12 .sum_lutc_input = "datac";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\R_src2_lo[11]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cycloneive_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[11]~q ),
	.cin(gnd),
	.combout(\Add1~29_combout ),
	.cout());
defparam \Add1~29 .lut_mask = 16'h0FF0;
defparam \Add1~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[10]~13 (
	.dataa(\D_iw[16]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[10]~13_combout ),
	.cout());
defparam \R_src2_lo[10]~13 .lut_mask = 16'hACFF;
defparam \R_src2_lo[10]~13 .sum_lutc_input = "datac";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\R_src2_lo[10]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cycloneive_lcell_comb \Add1~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[10]~q ),
	.cin(gnd),
	.combout(\Add1~30_combout ),
	.cout());
defparam \Add1~30 .lut_mask = 16'h0FF0;
defparam \Add1~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[9]~14 (
	.dataa(\D_iw[15]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[9]~14_combout ),
	.cout());
defparam \R_src2_lo[9]~14 .lut_mask = 16'hACFF;
defparam \R_src2_lo[9]~14 .sum_lutc_input = "datac";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\R_src2_lo[9]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cycloneive_lcell_comb \Add1~31 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[9]~q ),
	.cin(gnd),
	.combout(\Add1~31_combout ),
	.cout());
defparam \Add1~31 .lut_mask = 16'h0FF0;
defparam \Add1~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[8]~15 (
	.dataa(\D_iw[14]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[8]~15_combout ),
	.cout());
defparam \R_src2_lo[8]~15 .lut_mask = 16'hACFF;
defparam \R_src2_lo[8]~15 .sum_lutc_input = "datac";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\R_src2_lo[8]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cycloneive_lcell_comb \Add1~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[8]~q ),
	.cin(gnd),
	.combout(\Add1~32_combout ),
	.cout());
defparam \Add1~32 .lut_mask = 16'h0FF0;
defparam \Add1~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~33 (
	.dataa(\Add1~32_combout ),
	.datab(\E_src1[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~33_combout ),
	.cout(\Add1~34 ));
defparam \Add1~33 .lut_mask = 16'h967F;
defparam \Add1~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~35 (
	.dataa(\Add1~31_combout ),
	.datab(\E_src1[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~34 ),
	.combout(\Add1~35_combout ),
	.cout(\Add1~36 ));
defparam \Add1~35 .lut_mask = 16'h96EF;
defparam \Add1~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~37 (
	.dataa(\Add1~30_combout ),
	.datab(\E_src1[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~36 ),
	.combout(\Add1~37_combout ),
	.cout(\Add1~38 ));
defparam \Add1~37 .lut_mask = 16'h967F;
defparam \Add1~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~39 (
	.dataa(\Add1~29_combout ),
	.datab(\E_src1[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~38 ),
	.combout(\Add1~39_combout ),
	.cout(\Add1~40 ));
defparam \Add1~39 .lut_mask = 16'h96EF;
defparam \Add1~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~41 (
	.dataa(\Add1~28_combout ),
	.datab(\E_src1[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~40 ),
	.combout(\Add1~41_combout ),
	.cout(\Add1~42 ));
defparam \Add1~41 .lut_mask = 16'h967F;
defparam \Add1~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~43 (
	.dataa(\Add1~27_combout ),
	.datab(\E_src1[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~42 ),
	.combout(\Add1~43_combout ),
	.cout(\Add1~44 ));
defparam \Add1~43 .lut_mask = 16'h96EF;
defparam \Add1~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~45 (
	.dataa(\Add1~26_combout ),
	.datab(\E_src1[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~44 ),
	.combout(\Add1~45_combout ),
	.cout(\Add1~46 ));
defparam \Add1~45 .lut_mask = 16'h967F;
defparam \Add1~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[14]~1 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[14]~q ),
	.datac(\E_src1[14]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[14]~1_combout ),
	.cout());
defparam \E_logic_result[14]~1 .lut_mask = 16'h6996;
defparam \E_logic_result[14]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[14]~16 (
	.dataa(\Add1~45_combout ),
	.datab(\E_logic_result[14]~1_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[14]~16_combout ),
	.cout());
defparam \W_alu_result[14]~16 .lut_mask = 16'hAACC;
defparam \W_alu_result[14]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[13]~2 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[13]~q ),
	.datac(\E_src1[13]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[13]~2_combout ),
	.cout());
defparam \E_logic_result[13]~2 .lut_mask = 16'h6996;
defparam \E_logic_result[13]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[13]~17 (
	.dataa(\Add1~43_combout ),
	.datab(\E_logic_result[13]~2_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[13]~17_combout ),
	.cout());
defparam \W_alu_result[13]~17 .lut_mask = 16'hAACC;
defparam \W_alu_result[13]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[18]~10 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[18]~10_combout ),
	.cout());
defparam \E_src2[18]~10 .lut_mask = 16'hAACC;
defparam \E_src2[18]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~6_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~3 .lut_mask = 16'hFAFC;
defparam \D_ctrl_unsigned_lo_imm16~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~4 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_unsigned_lo_imm16~4 .sum_lutc_input = "datac";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cycloneive_lcell_comb \R_src2_hi~0 (
	.dataa(\R_ctrl_force_src2_zero~q ),
	.datab(\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_hi~0_combout ),
	.cout());
defparam \R_src2_hi~0 .lut_mask = 16'hEEEE;
defparam \R_src2_hi~0 .sum_lutc_input = "datac";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\E_src2[18]~10_combout ),
	.asdata(\D_iw[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cycloneive_lcell_comb \Add1~47 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[18]~q ),
	.cin(gnd),
	.combout(\Add1~47_combout ),
	.cout());
defparam \Add1~47 .lut_mask = 16'h0FF0;
defparam \Add1~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[17]~11 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[17]~11_combout ),
	.cout());
defparam \E_src2[17]~11 .lut_mask = 16'hAACC;
defparam \E_src2[17]~11 .sum_lutc_input = "datac";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\E_src2[17]~11_combout ),
	.asdata(\D_iw[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cycloneive_lcell_comb \Add1~48 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[17]~q ),
	.cin(gnd),
	.combout(\Add1~48_combout ),
	.cout());
defparam \Add1~48 .lut_mask = 16'h0FF0;
defparam \Add1~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[16]~12 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[16]~12_combout ),
	.cout());
defparam \E_src2[16]~12 .lut_mask = 16'hAACC;
defparam \E_src2[16]~12 .sum_lutc_input = "datac";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\E_src2[16]~12_combout ),
	.asdata(\D_iw[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cycloneive_lcell_comb \Add1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[16]~q ),
	.cin(gnd),
	.combout(\Add1~49_combout ),
	.cout());
defparam \Add1~49 .lut_mask = 16'h0FF0;
defparam \Add1~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[15]~16 (
	.dataa(\D_iw[21]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[12]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[15]~16_combout ),
	.cout());
defparam \R_src2_lo[15]~16 .lut_mask = 16'hACFF;
defparam \R_src2_lo[15]~16 .sum_lutc_input = "datac";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\R_src2_lo[15]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cycloneive_lcell_comb \Add1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[15]~q ),
	.cin(gnd),
	.combout(\Add1~50_combout ),
	.cout());
defparam \Add1~50 .lut_mask = 16'h0FF0;
defparam \Add1~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~51 (
	.dataa(\Add1~50_combout ),
	.datab(\E_src1[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~46 ),
	.combout(\Add1~51_combout ),
	.cout(\Add1~52 ));
defparam \Add1~51 .lut_mask = 16'h96EF;
defparam \Add1~51 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~53 (
	.dataa(\Add1~49_combout ),
	.datab(\E_src1[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~52 ),
	.combout(\Add1~53_combout ),
	.cout(\Add1~54 ));
defparam \Add1~53 .lut_mask = 16'h967F;
defparam \Add1~53 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~55 (
	.dataa(\Add1~48_combout ),
	.datab(\E_src1[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~54 ),
	.combout(\Add1~55_combout ),
	.cout(\Add1~56 ));
defparam \Add1~55 .lut_mask = 16'h96EF;
defparam \Add1~55 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~57 (
	.dataa(\Add1~47_combout ),
	.datab(\E_src1[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~56 ),
	.combout(\Add1~57_combout ),
	.cout(\Add1~58 ));
defparam \Add1~57 .lut_mask = 16'h967F;
defparam \Add1~57 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[18]~3 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[18]~q ),
	.datac(\E_src1[18]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[18]~3_combout ),
	.cout());
defparam \E_logic_result[18]~3 .lut_mask = 16'h6996;
defparam \E_logic_result[18]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[18]~12 (
	.dataa(\Add1~57_combout ),
	.datab(\E_logic_result[18]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[18]~12_combout ),
	.cout());
defparam \W_alu_result[18]~12 .lut_mask = 16'hAACC;
defparam \W_alu_result[18]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[17]~4 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[17]~q ),
	.datac(\E_src1[17]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[17]~4_combout ),
	.cout());
defparam \E_logic_result[17]~4 .lut_mask = 16'h6996;
defparam \E_logic_result[17]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[17]~13 (
	.dataa(\Add1~55_combout ),
	.datab(\E_logic_result[17]~4_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[17]~13_combout ),
	.cout());
defparam \W_alu_result[17]~13 .lut_mask = 16'hAACC;
defparam \W_alu_result[17]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[16]~5 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[16]~q ),
	.datac(\E_src1[16]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[16]~5_combout ),
	.cout());
defparam \E_logic_result[16]~5 .lut_mask = 16'h6996;
defparam \E_logic_result[16]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[16]~14 (
	.dataa(\Add1~53_combout ),
	.datab(\E_logic_result[16]~5_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[16]~14_combout ),
	.cout());
defparam \W_alu_result[16]~14 .lut_mask = 16'hAACC;
defparam \W_alu_result[16]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[15]~6 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[15]~q ),
	.datac(\E_src1[15]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[15]~6_combout ),
	.cout());
defparam \E_logic_result[15]~6 .lut_mask = 16'h6996;
defparam \E_logic_result[15]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[15]~15 (
	.dataa(\Add1~51_combout ),
	.datab(\E_logic_result[15]~6_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[15]~15_combout ),
	.cout());
defparam \W_alu_result[15]~15 .lut_mask = 16'hAACC;
defparam \W_alu_result[15]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[12]~7 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[12]~q ),
	.datac(\E_src1[12]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[12]~7_combout ),
	.cout());
defparam \E_logic_result[12]~7 .lut_mask = 16'h6996;
defparam \E_logic_result[12]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[12]~18 (
	.dataa(\Add1~41_combout ),
	.datab(\E_logic_result[12]~7_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[12]~18_combout ),
	.cout());
defparam \W_alu_result[12]~18 .lut_mask = 16'hAACC;
defparam \W_alu_result[12]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[11]~8 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[11]~q ),
	.datac(\E_src1[11]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[11]~8_combout ),
	.cout());
defparam \E_logic_result[11]~8 .lut_mask = 16'h6996;
defparam \E_logic_result[11]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[11]~19 (
	.dataa(\Add1~39_combout ),
	.datab(\E_logic_result[11]~8_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[11]~19_combout ),
	.cout());
defparam \W_alu_result[11]~19 .lut_mask = 16'hAACC;
defparam \W_alu_result[11]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[10]~9 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[10]~q ),
	.datac(\E_src1[10]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[10]~9_combout ),
	.cout());
defparam \E_logic_result[10]~9 .lut_mask = 16'h6996;
defparam \E_logic_result[10]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[10]~20 (
	.dataa(\Add1~37_combout ),
	.datab(\E_logic_result[10]~9_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[10]~20_combout ),
	.cout());
defparam \W_alu_result[10]~20 .lut_mask = 16'hAACC;
defparam \W_alu_result[10]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[9]~10 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[9]~q ),
	.datac(\E_src1[9]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[9]~10_combout ),
	.cout());
defparam \E_logic_result[9]~10 .lut_mask = 16'h6996;
defparam \E_logic_result[9]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[9]~21 (
	.dataa(\Add1~35_combout ),
	.datab(\E_logic_result[9]~10_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[9]~21_combout ),
	.cout());
defparam \W_alu_result[9]~21 .lut_mask = 16'hAACC;
defparam \W_alu_result[9]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[23]~5 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[23]~5_combout ),
	.cout());
defparam \E_src2[23]~5 .lut_mask = 16'hAACC;
defparam \E_src2[23]~5 .sum_lutc_input = "datac";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\E_src2[23]~5_combout ),
	.asdata(\D_iw[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cycloneive_lcell_comb \Add1~59 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[23]~q ),
	.cin(gnd),
	.combout(\Add1~59_combout ),
	.cout());
defparam \Add1~59 .lut_mask = 16'h0FF0;
defparam \Add1~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[22]~6 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[22]~6_combout ),
	.cout());
defparam \E_src2[22]~6 .lut_mask = 16'hAACC;
defparam \E_src2[22]~6 .sum_lutc_input = "datac";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\E_src2[22]~6_combout ),
	.asdata(\D_iw[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cycloneive_lcell_comb \Add1~60 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[22]~q ),
	.cin(gnd),
	.combout(\Add1~60_combout ),
	.cout());
defparam \Add1~60 .lut_mask = 16'h0FF0;
defparam \Add1~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[21]~7 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[21]~7_combout ),
	.cout());
defparam \E_src2[21]~7 .lut_mask = 16'hAACC;
defparam \E_src2[21]~7 .sum_lutc_input = "datac";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\E_src2[21]~7_combout ),
	.asdata(\D_iw[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cycloneive_lcell_comb \Add1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[21]~q ),
	.cin(gnd),
	.combout(\Add1~61_combout ),
	.cout());
defparam \Add1~61 .lut_mask = 16'h0FF0;
defparam \Add1~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[20]~8 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[20]~8_combout ),
	.cout());
defparam \E_src2[20]~8 .lut_mask = 16'hAACC;
defparam \E_src2[20]~8 .sum_lutc_input = "datac";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\E_src2[20]~8_combout ),
	.asdata(\D_iw[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cycloneive_lcell_comb \Add1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[20]~q ),
	.cin(gnd),
	.combout(\Add1~62_combout ),
	.cout());
defparam \Add1~62 .lut_mask = 16'h0FF0;
defparam \Add1~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[19]~9 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[19]~9_combout ),
	.cout());
defparam \E_src2[19]~9 .lut_mask = 16'hAACC;
defparam \E_src2[19]~9 .sum_lutc_input = "datac";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\E_src2[19]~9_combout ),
	.asdata(\D_iw[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cycloneive_lcell_comb \Add1~63 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[19]~q ),
	.cin(gnd),
	.combout(\Add1~63_combout ),
	.cout());
defparam \Add1~63 .lut_mask = 16'h0FF0;
defparam \Add1~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~64 (
	.dataa(\Add1~63_combout ),
	.datab(\E_src1[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~58 ),
	.combout(\Add1~64_combout ),
	.cout(\Add1~65 ));
defparam \Add1~64 .lut_mask = 16'h96EF;
defparam \Add1~64 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~66 (
	.dataa(\Add1~62_combout ),
	.datab(\E_src1[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~65 ),
	.combout(\Add1~66_combout ),
	.cout(\Add1~67 ));
defparam \Add1~66 .lut_mask = 16'h967F;
defparam \Add1~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~68 (
	.dataa(\Add1~61_combout ),
	.datab(\E_src1[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~67 ),
	.combout(\Add1~68_combout ),
	.cout(\Add1~69 ));
defparam \Add1~68 .lut_mask = 16'h96EF;
defparam \Add1~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~70 (
	.dataa(\Add1~60_combout ),
	.datab(\E_src1[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~69 ),
	.combout(\Add1~70_combout ),
	.cout(\Add1~71 ));
defparam \Add1~70 .lut_mask = 16'h967F;
defparam \Add1~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~72 (
	.dataa(\Add1~59_combout ),
	.datab(\E_src1[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~71 ),
	.combout(\Add1~72_combout ),
	.cout(\Add1~73 ));
defparam \Add1~72 .lut_mask = 16'h96EF;
defparam \Add1~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[23]~11 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[23]~q ),
	.datac(\E_src1[23]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[23]~11_combout ),
	.cout());
defparam \E_logic_result[23]~11 .lut_mask = 16'h6996;
defparam \E_logic_result[23]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[23]~5 (
	.dataa(\Add1~72_combout ),
	.datab(\E_logic_result[23]~11_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[23]~5_combout ),
	.cout());
defparam \W_alu_result[23]~5 .lut_mask = 16'hAACC;
defparam \W_alu_result[23]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[22]~12 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[22]~q ),
	.datac(\E_src1[22]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[22]~12_combout ),
	.cout());
defparam \E_logic_result[22]~12 .lut_mask = 16'h6996;
defparam \E_logic_result[22]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[22]~6 (
	.dataa(\Add1~70_combout ),
	.datab(\E_logic_result[22]~12_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[22]~6_combout ),
	.cout());
defparam \W_alu_result[22]~6 .lut_mask = 16'hAACC;
defparam \W_alu_result[22]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[8]~13 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[8]~q ),
	.datac(\E_src1[8]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[8]~13_combout ),
	.cout());
defparam \E_logic_result[8]~13 .lut_mask = 16'h6996;
defparam \E_logic_result[8]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[8]~22 (
	.dataa(\Add1~33_combout ),
	.datab(\E_logic_result[8]~13_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[8]~22_combout ),
	.cout());
defparam \W_alu_result[8]~22 .lut_mask = 16'hAACC;
defparam \W_alu_result[8]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[6]~14 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[6]~q ),
	.datac(\E_src1[6]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[6]~14_combout ),
	.cout());
defparam \E_logic_result[6]~14 .lut_mask = 16'h6996;
defparam \E_logic_result[6]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[6]~24 (
	.dataa(\Add1~22_combout ),
	.datab(\E_logic_result[6]~14_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[6]~24_combout ),
	.cout());
defparam \W_alu_result[6]~24 .lut_mask = 16'hAACC;
defparam \W_alu_result[6]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[24]~4 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[24]~4_combout ),
	.cout());
defparam \E_src2[24]~4 .lut_mask = 16'hAACC;
defparam \E_src2[24]~4 .sum_lutc_input = "datac";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\E_src2[24]~4_combout ),
	.asdata(\D_iw[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cycloneive_lcell_comb \Add1~74 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[24]~q ),
	.cin(gnd),
	.combout(\Add1~74_combout ),
	.cout());
defparam \Add1~74 .lut_mask = 16'h0FF0;
defparam \Add1~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~75 (
	.dataa(\Add1~74_combout ),
	.datab(\E_src1[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~73 ),
	.combout(\Add1~75_combout ),
	.cout(\Add1~76 ));
defparam \Add1~75 .lut_mask = 16'h967F;
defparam \Add1~75 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[24]~15 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[24]~q ),
	.datac(\E_src1[24]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[24]~15_combout ),
	.cout());
defparam \E_logic_result[24]~15 .lut_mask = 16'h6996;
defparam \E_logic_result[24]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[24]~4 (
	.dataa(\Add1~75_combout ),
	.datab(\E_logic_result[24]~15_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[24]~4_combout ),
	.cout());
defparam \W_alu_result[24]~4 .lut_mask = 16'hAACC;
defparam \W_alu_result[24]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[21]~16 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[21]~q ),
	.datac(\E_src1[21]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[21]~16_combout ),
	.cout());
defparam \E_logic_result[21]~16 .lut_mask = 16'h6996;
defparam \E_logic_result[21]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[21]~9 (
	.dataa(\Add1~68_combout ),
	.datab(\E_logic_result[21]~16_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[21]~9_combout ),
	.cout());
defparam \W_alu_result[21]~9 .lut_mask = 16'hAACC;
defparam \W_alu_result[21]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[20]~17 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[20]~q ),
	.datac(\E_src1[20]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[20]~17_combout ),
	.cout());
defparam \E_logic_result[20]~17 .lut_mask = 16'h6996;
defparam \E_logic_result[20]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[20]~10 (
	.dataa(\Add1~66_combout ),
	.datab(\E_logic_result[20]~17_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[20]~10_combout ),
	.cout());
defparam \W_alu_result[20]~10 .lut_mask = 16'hAACC;
defparam \W_alu_result[20]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[19]~18 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[19]~q ),
	.datac(\E_src1[19]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[19]~18_combout ),
	.cout());
defparam \E_logic_result[19]~18 .lut_mask = 16'h6996;
defparam \E_logic_result[19]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[19]~11 (
	.dataa(\Add1~64_combout ),
	.datab(\E_logic_result[19]~18_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[19]~11_combout ),
	.cout());
defparam \W_alu_result[19]~11 .lut_mask = 16'hAACC;
defparam \W_alu_result[19]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[28]~0 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[28]~0_combout ),
	.cout());
defparam \E_src2[28]~0 .lut_mask = 16'hAACC;
defparam \E_src2[28]~0 .sum_lutc_input = "datac";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\E_src2[28]~0_combout ),
	.asdata(\D_iw[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cycloneive_lcell_comb \Add1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[28]~q ),
	.cin(gnd),
	.combout(\Add1~77_combout ),
	.cout());
defparam \Add1~77 .lut_mask = 16'h0FF0;
defparam \Add1~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[27]~1 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[27]~1_combout ),
	.cout());
defparam \E_src2[27]~1 .lut_mask = 16'hAACC;
defparam \E_src2[27]~1 .sum_lutc_input = "datac";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\E_src2[27]~1_combout ),
	.asdata(\D_iw[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cycloneive_lcell_comb \Add1~78 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[27]~q ),
	.cin(gnd),
	.combout(\Add1~78_combout ),
	.cout());
defparam \Add1~78 .lut_mask = 16'h0FF0;
defparam \Add1~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[26]~2 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[26]~2_combout ),
	.cout());
defparam \E_src2[26]~2 .lut_mask = 16'hAACC;
defparam \E_src2[26]~2 .sum_lutc_input = "datac";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\E_src2[26]~2_combout ),
	.asdata(\D_iw[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cycloneive_lcell_comb \Add1~79 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[26]~q ),
	.cin(gnd),
	.combout(\Add1~79_combout ),
	.cout());
defparam \Add1~79 .lut_mask = 16'h0FF0;
defparam \Add1~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[25]~3 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[25]~3_combout ),
	.cout());
defparam \E_src2[25]~3 .lut_mask = 16'hAACC;
defparam \E_src2[25]~3 .sum_lutc_input = "datac";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\E_src2[25]~3_combout ),
	.asdata(\D_iw[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cycloneive_lcell_comb \Add1~80 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[25]~q ),
	.cin(gnd),
	.combout(\Add1~80_combout ),
	.cout());
defparam \Add1~80 .lut_mask = 16'h0FF0;
defparam \Add1~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~81 (
	.dataa(\Add1~80_combout ),
	.datab(\E_src1[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~76 ),
	.combout(\Add1~81_combout ),
	.cout(\Add1~82 ));
defparam \Add1~81 .lut_mask = 16'h96EF;
defparam \Add1~81 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~83 (
	.dataa(\Add1~79_combout ),
	.datab(\E_src1[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~82 ),
	.combout(\Add1~83_combout ),
	.cout(\Add1~84 ));
defparam \Add1~83 .lut_mask = 16'h967F;
defparam \Add1~83 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~85 (
	.dataa(\Add1~78_combout ),
	.datab(\E_src1[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~84 ),
	.combout(\Add1~85_combout ),
	.cout(\Add1~86 ));
defparam \Add1~85 .lut_mask = 16'h96EF;
defparam \Add1~85 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~87 (
	.dataa(\Add1~77_combout ),
	.datab(\E_src1[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~86 ),
	.combout(\Add1~87_combout ),
	.cout(\Add1~88 ));
defparam \Add1~87 .lut_mask = 16'h967F;
defparam \Add1~87 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[28]~19 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[28]~q ),
	.datac(\E_src1[28]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[28]~19_combout ),
	.cout());
defparam \E_logic_result[28]~19 .lut_mask = 16'h6996;
defparam \E_logic_result[28]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[28]~0 (
	.dataa(\Add1~87_combout ),
	.datab(\E_logic_result[28]~19_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[28]~0_combout ),
	.cout());
defparam \W_alu_result[28]~0 .lut_mask = 16'hAACC;
defparam \W_alu_result[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[27]~20 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[27]~q ),
	.datac(\E_src1[27]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[27]~20_combout ),
	.cout());
defparam \E_logic_result[27]~20 .lut_mask = 16'h6996;
defparam \E_logic_result[27]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[27]~1 (
	.dataa(\Add1~85_combout ),
	.datab(\E_logic_result[27]~20_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[27]~1_combout ),
	.cout());
defparam \W_alu_result[27]~1 .lut_mask = 16'hAACC;
defparam \W_alu_result[27]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[26]~21 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[26]~q ),
	.datac(\E_src1[26]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[26]~21_combout ),
	.cout());
defparam \E_logic_result[26]~21 .lut_mask = 16'h6996;
defparam \E_logic_result[26]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[26]~2 (
	.dataa(\Add1~83_combout ),
	.datab(\E_logic_result[26]~21_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[26]~2_combout ),
	.cout());
defparam \W_alu_result[26]~2 .lut_mask = 16'hAACC;
defparam \W_alu_result[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[25]~22 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[25]~q ),
	.datac(\E_src1[25]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[25]~22_combout ),
	.cout());
defparam \E_logic_result[25]~22 .lut_mask = 16'h6996;
defparam \E_logic_result[25]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[25]~3 (
	.dataa(\Add1~81_combout ),
	.datab(\E_logic_result[25]~22_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[25]~3_combout ),
	.cout());
defparam \W_alu_result[25]~3 .lut_mask = 16'hAACC;
defparam \W_alu_result[25]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[4]~23 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[4]~q ),
	.datac(\E_src1[4]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[4]~23_combout ),
	.cout());
defparam \E_logic_result[4]~23 .lut_mask = 16'h6996;
defparam \E_logic_result[4]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[4]~26 (
	.dataa(\Add1~18_combout ),
	.datab(\E_logic_result[4]~23_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[4]~26_combout ),
	.cout());
defparam \W_alu_result[4]~26 .lut_mask = 16'hAACC;
defparam \W_alu_result[4]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[5]~24 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[5]~q ),
	.datac(\E_src1[5]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[5]~24_combout ),
	.cout());
defparam \E_logic_result[5]~24 .lut_mask = 16'h6996;
defparam \E_logic_result[5]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[5]~25 (
	.dataa(\Add1~20_combout ),
	.datab(\E_logic_result[5]~24_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[5]~25_combout ),
	.cout());
defparam \W_alu_result[5]~25 .lut_mask = 16'hAACC;
defparam \W_alu_result[5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[2]~25 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[2]~q ),
	.datac(\E_src1[2]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[2]~25_combout ),
	.cout());
defparam \E_logic_result[2]~25 .lut_mask = 16'h6996;
defparam \E_logic_result[2]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[2]~7 (
	.dataa(\Add1~14_combout ),
	.datab(\E_logic_result[2]~25_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[2]~7_combout ),
	.cout());
defparam \W_alu_result[2]~7 .lut_mask = 16'hAACC;
defparam \W_alu_result[2]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[3]~26 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[3]~q ),
	.datac(\E_src1[3]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[3]~26_combout ),
	.cout());
defparam \E_logic_result[3]~26 .lut_mask = 16'h6996;
defparam \E_logic_result[3]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[3]~8 (
	.dataa(\Add1~16_combout ),
	.datab(\E_logic_result[3]~26_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[3]~8_combout ),
	.cout());
defparam \W_alu_result[3]~8 .lut_mask = 16'hAACC;
defparam \W_alu_result[3]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[24]~0 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[24]~0_combout ),
	.cout());
defparam \d_writedata[24]~0 .lut_mask = 16'hAACC;
defparam \d_writedata[24]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.cout());
defparam \D_ctrl_mem8~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~1 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.cout());
defparam \D_ctrl_mem8~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[25]~1 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[25]~1_combout ),
	.cout());
defparam \d_writedata[25]~1 .lut_mask = 16'hAACC;
defparam \d_writedata[25]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[26]~2 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[26]~2_combout ),
	.cout());
defparam \d_writedata[26]~2 .lut_mask = 16'hAACC;
defparam \d_writedata[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[27]~3 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[27]~3_combout ),
	.cout());
defparam \d_writedata[27]~3 .lut_mask = 16'hAACC;
defparam \d_writedata[27]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[28]~4 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[28]~4_combout ),
	.cout());
defparam \d_writedata[28]~4 .lut_mask = 16'hAACC;
defparam \d_writedata[28]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[29]~5 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[29]~5_combout ),
	.cout());
defparam \d_writedata[29]~5 .lut_mask = 16'hAACC;
defparam \d_writedata[29]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[30]~6 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[30]~6_combout ),
	.cout());
defparam \d_writedata[30]~6 .lut_mask = 16'hAACC;
defparam \d_writedata[30]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[31]~7 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[31]~7_combout ),
	.cout());
defparam \d_writedata[31]~7 .lut_mask = 16'hAACC;
defparam \d_writedata[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb E_st_stall(
	.dataa(d_write1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_st~q ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\E_st_stall~combout ),
	.cout());
defparam E_st_stall.lut_mask = 16'hFFFE;
defparam E_st_stall.sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[8]~0 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[8]~0_combout ),
	.cout());
defparam \E_st_data[8]~0 .lut_mask = 16'hEFFE;
defparam \E_st_data[8]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[9]~1 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[9]~1_combout ),
	.cout());
defparam \E_st_data[9]~1 .lut_mask = 16'hEFFE;
defparam \E_st_data[9]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[10]~2 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[10]~2_combout ),
	.cout());
defparam \E_st_data[10]~2 .lut_mask = 16'hEFFE;
defparam \E_st_data[10]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[11]~3 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[11]~3_combout ),
	.cout());
defparam \E_st_data[11]~3 .lut_mask = 16'hEFFE;
defparam \E_st_data[11]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[12]~4 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[12]~4_combout ),
	.cout());
defparam \E_st_data[12]~4 .lut_mask = 16'hEFFE;
defparam \E_st_data[12]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[13]~5 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[13]~5_combout ),
	.cout());
defparam \E_st_data[13]~5 .lut_mask = 16'hEFFE;
defparam \E_st_data[13]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[14]~6 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[14]~6_combout ),
	.cout());
defparam \E_st_data[14]~6 .lut_mask = 16'hEFFE;
defparam \E_st_data[14]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[15]~7 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[15]~7_combout ),
	.cout());
defparam \E_st_data[15]~7 .lut_mask = 16'hEFFE;
defparam \E_st_data[15]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[23]~8 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(\D_ctrl_mem16~0_combout ),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\d_writedata[23]~8_combout ),
	.cout());
defparam \d_writedata[23]~8 .lut_mask = 16'hEEFF;
defparam \d_writedata[23]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[16]~8 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[16]~8_combout ),
	.cout());
defparam \E_st_data[16]~8 .lut_mask = 16'hAACC;
defparam \E_st_data[16]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[17]~9 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[17]~9_combout ),
	.cout());
defparam \E_st_data[17]~9 .lut_mask = 16'hAACC;
defparam \E_st_data[17]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_read_nxt~0 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(d_read1),
	.datad(av_ld_getting_data),
	.cin(gnd),
	.combout(\d_read_nxt~0_combout ),
	.cout());
defparam \d_read_nxt~0 .lut_mask = 16'hFEFF;
defparam \d_read_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_uncond_cti_non_br~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~2 (
	.dataa(\D_ctrl_jmp_direct~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~1_combout ),
	.datac(gnd),
	.datad(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~2_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~2 .lut_mask = 16'hEEFF;
defparam \D_ctrl_uncond_cti_non_br~2 .sum_lutc_input = "datac";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(clk_clk),
	.d(\D_ctrl_uncond_cti_non_br~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cycloneive_lcell_comb \Equal0~20 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~20_combout ),
	.cout());
defparam \Equal0~20 .lut_mask = 16'hF7F7;
defparam \Equal0~20 .sum_lutc_input = "datac";

dffeas R_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\Equal0~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

dffeas \R_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.cout());
defparam \D_logic_op_raw[0]~1 .lut_mask = 16'hEFFE;
defparam \D_logic_op_raw[0]~1 .sum_lutc_input = "datac";

dffeas \R_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cycloneive_lcell_comb \Equal127~0 (
	.dataa(\E_logic_result[28]~19_combout ),
	.datab(\E_logic_result[27]~20_combout ),
	.datac(\E_logic_result[26]~21_combout ),
	.datad(\E_logic_result[25]~22_combout ),
	.cin(gnd),
	.combout(\Equal127~0_combout ),
	.cout());
defparam \Equal127~0 .lut_mask = 16'h7FFF;
defparam \Equal127~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~1 (
	.dataa(\E_logic_result[23]~11_combout ),
	.datab(\E_logic_result[22]~12_combout ),
	.datac(\E_logic_result[24]~15_combout ),
	.datad(\E_logic_result[21]~16_combout ),
	.cin(gnd),
	.combout(\Equal127~1_combout ),
	.cout());
defparam \Equal127~1 .lut_mask = 16'h7FFF;
defparam \Equal127~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~2 (
	.dataa(\E_logic_result[20]~17_combout ),
	.datab(\E_logic_result[19]~18_combout ),
	.datac(\E_logic_result[18]~3_combout ),
	.datad(\E_logic_result[17]~4_combout ),
	.cin(gnd),
	.combout(\Equal127~2_combout ),
	.cout());
defparam \Equal127~2 .lut_mask = 16'h7FFF;
defparam \Equal127~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~3 (
	.dataa(\E_logic_result[14]~1_combout ),
	.datab(\E_logic_result[13]~2_combout ),
	.datac(\E_logic_result[16]~5_combout ),
	.datad(\E_logic_result[15]~6_combout ),
	.cin(gnd),
	.combout(\Equal127~3_combout ),
	.cout());
defparam \Equal127~3 .lut_mask = 16'h7FFF;
defparam \Equal127~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~4 (
	.dataa(\Equal127~0_combout ),
	.datab(\Equal127~1_combout ),
	.datac(\Equal127~2_combout ),
	.datad(\Equal127~3_combout ),
	.cin(gnd),
	.combout(\Equal127~4_combout ),
	.cout());
defparam \Equal127~4 .lut_mask = 16'hFFFE;
defparam \Equal127~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~5 (
	.dataa(\E_logic_result[12]~7_combout ),
	.datab(\E_logic_result[11]~8_combout ),
	.datac(\E_logic_result[10]~9_combout ),
	.datad(\E_logic_result[9]~10_combout ),
	.cin(gnd),
	.combout(\Equal127~5_combout ),
	.cout());
defparam \Equal127~5 .lut_mask = 16'h7FFF;
defparam \Equal127~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~6 (
	.dataa(\E_logic_result[5]~24_combout ),
	.datab(\E_logic_result[7]~0_combout ),
	.datac(\E_logic_result[8]~13_combout ),
	.datad(\E_logic_result[6]~14_combout ),
	.cin(gnd),
	.combout(\Equal127~6_combout ),
	.cout());
defparam \Equal127~6 .lut_mask = 16'h7FFF;
defparam \Equal127~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[0]~27 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[0]~q ),
	.datac(\E_src1[0]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[0]~27_combout ),
	.cout());
defparam \E_logic_result[0]~27 .lut_mask = 16'h6996;
defparam \E_logic_result[0]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~7 (
	.dataa(\E_logic_result[4]~23_combout ),
	.datab(\E_logic_result[2]~25_combout ),
	.datac(\E_logic_result[3]~26_combout ),
	.datad(\E_logic_result[0]~27_combout ),
	.cin(gnd),
	.combout(\Equal127~7_combout ),
	.cout());
defparam \Equal127~7 .lut_mask = 16'h7FFF;
defparam \Equal127~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~1 (
	.dataa(\D_iw[21]~q ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\R_ctrl_hi_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~1_combout ),
	.cout());
defparam \R_src2_hi[15]~1 .lut_mask = 16'hEFFE;
defparam \R_src2_hi[15]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~2 (
	.dataa(\R_src2_hi[15]~1_combout ),
	.datab(gnd),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(\R_ctrl_unsigned_lo_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~2_combout ),
	.cout());
defparam \R_src2_hi[15]~2 .lut_mask = 16'hAFFF;
defparam \R_src2_hi[15]~2 .sum_lutc_input = "datac";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\R_src2_hi[15]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[31]~28 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_src1[31]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[31]~28_combout ),
	.cout());
defparam \E_logic_result[31]~28 .lut_mask = 16'h6996;
defparam \E_logic_result[31]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[29]~13 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[29]~13_combout ),
	.cout());
defparam \E_src2[29]~13 .lut_mask = 16'hAACC;
defparam \E_src2[29]~13 .sum_lutc_input = "datac";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\E_src2[29]~13_combout ),
	.asdata(\D_iw[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[29]~29 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[29]~q ),
	.datac(\E_src1[29]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[29]~29_combout ),
	.cout());
defparam \E_logic_result[29]~29 .lut_mask = 16'h6996;
defparam \E_logic_result[29]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[1]~30 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[1]~q ),
	.datac(\E_src1[1]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[1]~30_combout ),
	.cout());
defparam \E_logic_result[1]~30 .lut_mask = 16'h6996;
defparam \E_logic_result[1]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[30]~14 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[30]~14_combout ),
	.cout());
defparam \E_src2[30]~14 .lut_mask = 16'hAACC;
defparam \E_src2[30]~14 .sum_lutc_input = "datac";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\E_src2[30]~14_combout ),
	.asdata(\D_iw[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[30]~31 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[30]~q ),
	.datac(\E_src1[30]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[30]~31_combout ),
	.cout());
defparam \E_logic_result[30]~31 .lut_mask = 16'h6996;
defparam \E_logic_result[30]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~8 (
	.dataa(\E_logic_result[31]~28_combout ),
	.datab(\E_logic_result[29]~29_combout ),
	.datac(\E_logic_result[1]~30_combout ),
	.datad(\E_logic_result[30]~31_combout ),
	.cin(gnd),
	.combout(\Equal127~8_combout ),
	.cout());
defparam \Equal127~8 .lut_mask = 16'h7FFF;
defparam \Equal127~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~9 (
	.dataa(\Equal127~5_combout ),
	.datab(\Equal127~6_combout ),
	.datac(\Equal127~7_combout ),
	.datad(\Equal127~8_combout ),
	.cin(gnd),
	.combout(\Equal127~9_combout ),
	.cout());
defparam \Equal127~9 .lut_mask = 16'hFFFE;
defparam \Equal127~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_cmp_result~0 (
	.dataa(\R_compare_op[1]~q ),
	.datab(\R_compare_op[0]~q ),
	.datac(\Equal127~4_combout ),
	.datad(\Equal127~9_combout ),
	.cin(gnd),
	.combout(\E_cmp_result~0_combout ),
	.cout());
defparam \E_cmp_result~0 .lut_mask = 16'h6996;
defparam \E_cmp_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.cout());
defparam \E_invert_arith_src_msb~0 .lut_mask = 16'hEFFE;
defparam \E_invert_arith_src_msb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(\R_valid~q ),
	.datab(\E_invert_arith_src_msb~0_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_alu_subtract~8_combout ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.cout());
defparam \E_invert_arith_src_msb~1 .lut_mask = 16'hEFFF;
defparam \E_invert_arith_src_msb~1 .sum_lutc_input = "datac";

dffeas E_invert_arith_src_msb(
	.clk(clk_clk),
	.d(\E_invert_arith_src_msb~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cycloneive_lcell_comb \Add1~89 (
	.dataa(\E_alu_sub~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add1~89_combout ),
	.cout());
defparam \Add1~89 .lut_mask = 16'h9696;
defparam \Add1~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_arith_src1[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(\E_src1[31]~q ),
	.cin(gnd),
	.combout(\E_arith_src1[31]~combout ),
	.cout());
defparam \E_arith_src1[31] .lut_mask = 16'h0FF0;
defparam \E_arith_src1[31] .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~90 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[30]~q ),
	.cin(gnd),
	.combout(\Add1~90_combout ),
	.cout());
defparam \Add1~90 .lut_mask = 16'h0FF0;
defparam \Add1~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~91 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[29]~q ),
	.cin(gnd),
	.combout(\Add1~91_combout ),
	.cout());
defparam \Add1~91 .lut_mask = 16'h0FF0;
defparam \Add1~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~98 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~97 ),
	.combout(\Add1~98_combout ),
	.cout());
defparam \Add1~98 .lut_mask = 16'h5A5A;
defparam \Add1~98 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_cmp_result~1 (
	.dataa(\E_cmp_result~0_combout ),
	.datab(\R_compare_op[1]~q ),
	.datac(\Add1~98_combout ),
	.datad(\R_compare_op[0]~q ),
	.cin(gnd),
	.combout(\E_cmp_result~1_combout ),
	.cout());
defparam \E_cmp_result~1 .lut_mask = 16'hEBBE;
defparam \E_cmp_result~1 .sum_lutc_input = "datac";

dffeas W_cmp_result(
	.clk(clk_clk),
	.d(\E_cmp_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cycloneive_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(\R_ctrl_uncond_cti_non_br~q ),
	.datab(\R_ctrl_br_uncond~q ),
	.datac(\W_cmp_result~q ),
	.datad(\R_ctrl_br~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.cout());
defparam \F_pc_sel_nxt~0 .lut_mask = 16'hFFFE;
defparam \F_pc_sel_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[26]~6 (
	.dataa(\R_ctrl_break~q ),
	.datab(\F_pc_plus_one[26]~52_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[26]~6_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[26]~6 .lut_mask = 16'hEFFF;
defparam \F_pc_no_crst_nxt[26]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[26]~7 (
	.dataa(\F_pc_no_crst_nxt[26]~6_combout ),
	.datab(\Add1~87_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[26]~7_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[26]~7 .lut_mask = 16'hFEFF;
defparam \F_pc_no_crst_nxt[26]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[25]~34 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\R_ctrl_break~q ),
	.datad(\F_pc_plus_one[25]~50_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[25]~34_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[25]~34 .lut_mask = 16'hFFDF;
defparam \F_pc_no_crst_nxt[25]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(gnd),
	.datac(\R_ctrl_exception~q ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~0 .lut_mask = 16'hAFFF;
defparam \F_pc_sel_nxt.10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[25]~8 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\F_pc_no_crst_nxt[25]~34_combout ),
	.datac(\Add1~85_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[25]~8_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[25]~8 .lut_mask = 16'h7FFF;
defparam \F_pc_no_crst_nxt[25]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[24]~9 (
	.dataa(\Add1~83_combout ),
	.datab(\F_pc_plus_one[24]~48_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[24]~9_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[24]~9 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[24]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[23]~10 (
	.dataa(\Add1~81_combout ),
	.datab(\F_pc_plus_one[23]~46_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[23]~10_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[23]~10 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[23]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[22]~35 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\R_ctrl_break~q ),
	.datad(\F_pc_plus_one[22]~44_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[22]~35_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[22]~35 .lut_mask = 16'hFFFB;
defparam \F_pc_no_crst_nxt[22]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[22]~11 (
	.dataa(\R_ctrl_break~q ),
	.datab(\Add1~75_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_no_crst_nxt[22]~35_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[22]~11_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[22]~11 .lut_mask = 16'hFFEF;
defparam \F_pc_no_crst_nxt[22]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[21]~12 (
	.dataa(\Add1~72_combout ),
	.datab(\F_pc_plus_one[21]~42_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[21]~12_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[21]~12 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[21]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[20]~13 (
	.dataa(\Add1~70_combout ),
	.datab(\F_pc_plus_one[20]~40_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[20]~13_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[20]~13 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[20]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[19]~14 (
	.dataa(\Add1~68_combout ),
	.datab(\F_pc_plus_one[19]~38_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[19]~14_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[19]~14 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[19]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[18]~15 (
	.dataa(\Add1~66_combout ),
	.datab(\F_pc_plus_one[18]~36_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[18]~15_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[18]~15 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[18]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[17]~16 (
	.dataa(\Add1~64_combout ),
	.datab(\F_pc_plus_one[17]~34_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[17]~16_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[17]~16 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[17]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[16]~17 (
	.dataa(\Add1~57_combout ),
	.datab(\F_pc_plus_one[16]~32_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[16]~17_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[16]~17 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[16]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[15]~18 (
	.dataa(\Add1~55_combout ),
	.datab(\F_pc_plus_one[15]~30_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[15]~18_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[15]~18 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[15]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[14]~19 (
	.dataa(\Add1~53_combout ),
	.datab(\F_pc_plus_one[14]~28_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[14]~19_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[14]~19 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[14]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[13]~20 (
	.dataa(\Add1~51_combout ),
	.datab(\F_pc_plus_one[13]~26_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~20_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~20 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[13]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[12]~21 (
	.dataa(\Add1~45_combout ),
	.datab(\F_pc_plus_one[12]~24_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[12]~21_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[12]~21 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[12]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[11]~22 (
	.dataa(\Add1~43_combout ),
	.datab(\F_pc_plus_one[11]~22_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[11]~22_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[11]~22 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[11]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[10]~23 (
	.dataa(\Add1~41_combout ),
	.datab(\F_pc_plus_one[10]~20_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~23_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~23 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[10]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~36 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\R_ctrl_break~q ),
	.datad(\F_pc_plus_one[9]~18_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~36_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~36 .lut_mask = 16'hFFFD;
defparam \F_pc_no_crst_nxt[9]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~24 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\Add1~39_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_no_crst_nxt[9]~36_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~24_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~24 .lut_mask = 16'hFFFD;
defparam \F_pc_no_crst_nxt[9]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[8]~25 (
	.dataa(\Add1~37_combout ),
	.datab(\F_pc_plus_one[8]~16_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[8]~25_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[8]~25 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[8]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[7]~26 (
	.dataa(\Add1~35_combout ),
	.datab(\F_pc_plus_one[7]~14_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[7]~26_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[7]~26 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[7]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[5]~27 (
	.dataa(\Add1~24_combout ),
	.datab(\F_pc_plus_one[5]~10_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[5]~27_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[5]~27 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[5]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[6]~28 (
	.dataa(\Add1~33_combout ),
	.datab(\F_pc_plus_one[6]~12_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[6]~28_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[6]~28 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[6]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[4]~29 (
	.dataa(\Add1~22_combout ),
	.datab(\F_pc_plus_one[4]~8_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[4]~29_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[4]~29 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[4]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[1]~30 (
	.dataa(\Add1~16_combout ),
	.datab(\F_pc_plus_one[1]~2_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[1]~30_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[1]~30 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[1]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[3]~31 (
	.dataa(\F_pc_sel_nxt.10~1_combout ),
	.datab(\Add1~20_combout ),
	.datac(\F_pc_plus_one[3]~6_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[3]~31_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[3]~31 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[3]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_read_nxt~0 (
	.dataa(\W_valid~q ),
	.datab(gnd),
	.datac(i_read1),
	.datad(av_readdatavalid2),
	.cin(gnd),
	.combout(\i_read_nxt~0_combout ),
	.cout());
defparam \i_read_nxt~0 .lut_mask = 16'hFFF5;
defparam \i_read_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[2]~32 (
	.dataa(\Add1~18_combout ),
	.datab(\F_pc_plus_one[2]~4_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[2]~32_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[2]~32 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[2]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[0]~33 (
	.dataa(\Add1~14_combout ),
	.datab(\F_pc_plus_one[0]~0_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_sel_nxt.10~1_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[0]~33_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[0]~33 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[0]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \hbreak_enabled~0 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~10_combout ),
	.datac(hbreak_enabled1),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.cout());
defparam \hbreak_enabled~0 .lut_mask = 16'hFFF7;
defparam \hbreak_enabled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[0]~0 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~10_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[0]~0_combout ),
	.cout());
defparam \E_mem_byte_en[0]~0 .lut_mask = 16'h6FFF;
defparam \E_mem_byte_en[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[1]~1 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~10_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[1]~1_combout ),
	.cout());
defparam \E_mem_byte_en[1]~1 .lut_mask = 16'hF6FF;
defparam \E_mem_byte_en[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[2]~2 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~12_combout ),
	.datac(\D_ctrl_mem8~1_combout ),
	.datad(\Add1~10_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[2]~2_combout ),
	.cout());
defparam \E_mem_byte_en[2]~2 .lut_mask = 16'hDEFF;
defparam \E_mem_byte_en[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~12_combout ),
	.datac(\Add1~10_combout ),
	.datad(\D_ctrl_mem8~1_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.cout());
defparam \E_mem_byte_en[3]~3 .lut_mask = 16'hFDFE;
defparam \E_mem_byte_en[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[18]~10 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[18]~10_combout ),
	.cout());
defparam \E_st_data[18]~10 .lut_mask = 16'hAACC;
defparam \E_st_data[18]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[19]~11 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[19]~11_combout ),
	.cout());
defparam \E_st_data[19]~11 .lut_mask = 16'hAACC;
defparam \E_st_data[19]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[20]~12 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[20]~12_combout ),
	.cout());
defparam \E_st_data[20]~12 .lut_mask = 16'hAACC;
defparam \E_st_data[20]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[21]~13 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[21]~13_combout ),
	.cout());
defparam \E_st_data[21]~13 .lut_mask = 16'hAACC;
defparam \E_st_data[21]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[22]~14 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[22]~14_combout ),
	.cout());
defparam \E_st_data[22]~14 .lut_mask = 16'hAACC;
defparam \E_st_data[22]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[23]~15 (
	.dataa(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(\usb_system_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\d_writedata[23]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[23]~15_combout ),
	.cout());
defparam \E_st_data[23]~15 .lut_mask = 16'hAACC;
defparam \E_st_data[23]~15 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_cpu_cpu_nios2_oci (
	sr_0,
	jtag_break,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_5,
	readdata_6,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	resetrequest,
	waitrequest,
	mem_used_1,
	WideOr1,
	local_read,
	hbreak_enabled,
	mem,
	address_nxt,
	oci_ienable_6,
	oci_ienable_5,
	oci_single_step_mode,
	readdata_4,
	r_early_rst,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_14,
	readdata_15,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_20,
	readdata_18,
	readdata_19,
	readdata_17,
	readdata_21,
	readdata_27,
	readdata_28,
	readdata_31,
	readdata_30,
	readdata_29,
	debugaccess_nxt,
	writedata_nxt,
	byteenable_nxt,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	jtag_break;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_5;
output 	readdata_6;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
output 	resetrequest;
output 	waitrequest;
input 	mem_used_1;
input 	WideOr1;
input 	local_read;
input 	hbreak_enabled;
input 	mem;
input 	[8:0] address_nxt;
output 	oci_ienable_6;
output 	oci_ienable_5;
output 	oci_single_step_mode;
output 	readdata_4;
input 	r_early_rst;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_14;
output 	readdata_15;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_20;
output 	readdata_18;
output 	readdata_19;
output 	readdata_17;
output 	readdata_21;
output 	readdata_27;
output 	readdata_28;
output 	readdata_31;
output 	readdata_30;
output 	readdata_29;
input 	debugaccess_nxt;
input 	[31:0] writedata_nxt;
input 	[3:0] byteenable_nxt;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_no_action_break_a~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_usb_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ;
wire \write~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \read~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \debugaccess~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|ociram_wr_en~0_combout ;
wire \writedata[0]~q ;
wire \address[1]~q ;
wire \address[2]~q ;
wire \address[3]~q ;
wire \address[4]~q ;
wire \address[5]~q ;
wire \address[6]~q ;
wire \address[7]~q ;
wire \byteenable[0]~q ;
wire \the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ;
wire \the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ;
wire \the_usb_system_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \writedata[6]~q ;
wire \writedata[5]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \writedata[3]~q ;
wire \the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[22]~q ;
wire \the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ;
wire \the_usb_system_cpu_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \writedata[1]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \writedata[2]~q ;
wire \writedata[4]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \writedata[21]~q ;
wire \byteenable[2]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \writedata[22]~q ;
wire \writedata[23]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \writedata[25]~q ;
wire \writedata[26]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \writedata[13]~q ;
wire \writedata[16]~q ;
wire \writedata[12]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \writedata[14]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \writedata[10]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \writedata[9]~q ;
wire \writedata[8]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \writedata[7]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \writedata[20]~q ;
wire \writedata[18]~q ;
wire \writedata[19]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \writedata[17]~q ;
wire \writedata[27]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \writedata[28]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \writedata[31]~q ;
wire \the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \writedata[30]~q ;
wire \writedata[29]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \address[0]~q ;
wire \readdata~0_combout ;
wire \readdata~1_combout ;
wire \address[8]~q ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~15_combout ;
wire \readdata~22_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \readdata~8_combout ;
wire \readdata~9_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~16_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;
wire \readdata~20_combout ;
wire \readdata~21_combout ;
wire \readdata~23_combout ;
wire \readdata~24_combout ;
wire \readdata~25_combout ;
wire \readdata~26_combout ;
wire \readdata~27_combout ;
wire \readdata~28_combout ;
wire \readdata~29_combout ;
wire \readdata~30_combout ;
wire \readdata~31_combout ;
wire \readdata~32_combout ;


usb_system_usb_system_cpu_cpu_debug_slave_wrapper the_usb_system_cpu_cpu_debug_slave_wrapper(
	.sr_0(sr_0),
	.MonDReg_0(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.MonDReg_2(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.MonDReg_3(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.MonDReg_4(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_27(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_11(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_10(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_8(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_29(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.jdo_22(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_35(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_34(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.break_readreg_0(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.hbreak_enabled(hbreak_enabled),
	.break_readreg_1(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_37(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.jdo_36(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.take_no_action_break_a(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_no_action_break_a~0_combout ),
	.jdo_3(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.take_action_ocimem_b(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.monitor_ready(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_17(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.break_readreg_21(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.MonDReg_21(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.monitor_error(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.break_readreg_2(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_33(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_19(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_22(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.MonDReg_22(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.jdo_24(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_3(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.break_readreg_16(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_20(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.jdo_23(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_23(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.MonDReg_23(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.break_readreg_4(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_27(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_24(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_13(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_15(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_9(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_7(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_17(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_28(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_31(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_30(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_17(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.resetlatch(\the_usb_system_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.break_readreg_31(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_30(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_29(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_18(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.jdo_7(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.break_readreg_5(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_14(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_6(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_nios2_ocimem the_usb_system_cpu_cpu_nios2_ocimem(
	.MonDReg_0(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.q_a_0(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.MonDReg_2(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.q_a_1(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_21(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.MonDReg_3(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.q_a_22(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_11(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_5(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_10(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_20(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_18(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_19(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_17(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_27(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_31(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_30(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_29(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.MonDReg_4(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_27(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_11(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_10(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_8(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_29(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.waitrequest1(waitrequest),
	.jdo_22(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_35(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_34(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.MonDReg_1(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.take_action_ocimem_b(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.jdo_17(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.MonDReg_21(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.jdo_4(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.debugaccess(\debugaccess~q ),
	.ociram_wr_en(\the_usb_system_cpu_cpu_nios2_ocimem|ociram_wr_en~0_combout ),
	.r_early_rst(r_early_rst),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_25(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_33(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_5(\writedata[5]~q ),
	.jdo_19(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.writedata_3(\writedata[3]~q ),
	.MonDReg_22(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.jdo_24(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_5(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.MonDReg_16(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_20(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.jdo_23(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.writedata_2(\writedata[2]~q ),
	.writedata_4(\writedata[4]~q ),
	.MonDReg_23(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.writedata_21(\writedata[21]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.jdo_6(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.MonDReg_25(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_26(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_24(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.writedata_22(\writedata[22]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.MonDReg_13(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_16(\writedata[16]~q ),
	.writedata_12(\writedata[12]~q ),
	.MonDReg_14(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.writedata_14(\writedata[14]~q ),
	.MonDReg_15(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_10(\writedata[10]~q ),
	.MonDReg_9(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_8(\writedata[8]~q ),
	.MonDReg_7(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.writedata_7(\writedata[7]~q ),
	.MonDReg_6(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_19(\writedata[19]~q ),
	.MonDReg_17(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.writedata_17(\writedata[17]~q ),
	.writedata_27(\writedata[27]~q ),
	.MonDReg_28(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.writedata_28(\writedata[28]~q ),
	.MonDReg_31(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.writedata_31(\writedata[31]~q ),
	.MonDReg_30(\the_usb_system_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_29(\writedata[29]~q ),
	.jdo_16(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.jdo_7(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_14(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_nios2_avalon_reg the_usb_system_cpu_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.address_8(\address[8]~q ),
	.oci_ienable_6(oci_ienable_6),
	.oci_ienable_5(oci_ienable_5),
	.oci_single_step_mode1(oci_single_step_mode),
	.ociram_wr_en(\the_usb_system_cpu_cpu_nios2_ocimem|ociram_wr_en~0_combout ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.Equal0(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.Equal01(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.take_action_ocireg(\the_usb_system_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.writedata_6(\writedata[6]~q ),
	.writedata_5(\writedata[5]~q ),
	.writedata_3(\writedata[3]~q ),
	.oci_ienable_22(\the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[22]~q ),
	.Equal02(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_nios2_oci_break the_usb_system_cpu_cpu_nios2_oci_break(
	.jdo_22(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.break_readreg_0(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.jdo_0(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_37(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.jdo_36(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.take_no_action_break_a(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_no_action_break_a~0_combout ),
	.jdo_3(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_17(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.break_readreg_21(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_2(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_31(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_19(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_22(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.jdo_24(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_3(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.break_readreg_16(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_20(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.jdo_23(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_23(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_4(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_24(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_17(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.break_readreg_31(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_30(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_29(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_18(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.jdo_7(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.break_readreg_5(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_14(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_6(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_usb_system_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_nios2_oci_debug the_usb_system_cpu_cpu_nios2_oci_debug(
	.jtag_break1(jtag_break),
	.r_sync_rst(r_sync_rst),
	.resetrequest1(resetrequest),
	.jdo_22(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_35(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_34(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.monitor_ready1(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_21(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.monitor_error1(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_usb_system_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_25(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_19(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_go1(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.jdo_24(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_23(\the_usb_system_cpu_cpu_debug_slave_wrapper|the_usb_system_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.resetlatch1(\the_usb_system_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(waitrequest),
	.datab(WideOr1),
	.datac(mem),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFAFC;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(waitrequest),
	.datab(\read~q ),
	.datac(local_read),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hB8FF;
defparam \read~0 .sum_lutc_input = "datac";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~4_combout ),
	.asdata(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\readdata~15_combout ),
	.asdata(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\readdata~22_combout ),
	.asdata(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\readdata~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\readdata~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\readdata~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\readdata~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\readdata~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\readdata~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\readdata~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\readdata~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\readdata~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\readdata~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\readdata~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\address[0]~q ),
	.datab(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.datac(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datad(\the_usb_system_cpu_cpu_nios2_avalon_reg|oci_ienable[22]~q ),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hFFFE;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~1 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.datac(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hFEFE;
defparam \readdata~1 .sum_lutc_input = "datac";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.datac(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hFEFE;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(\the_usb_system_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hFEFE;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\readdata~0_combout ),
	.datab(oci_single_step_mode),
	.datac(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hFEFE;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\address[0]~q ),
	.datab(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.datac(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datad(oci_ienable_5),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hFEFF;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~22 (
	.dataa(\address[0]~q ),
	.datab(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~0_combout ),
	.datac(\the_usb_system_cpu_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datad(oci_ienable_6),
	.cin(gnd),
	.combout(\readdata~22_combout ),
	.cout());
defparam \readdata~22 .lut_mask = 16'hFEFF;
defparam \readdata~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hAACC;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hAACC;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hAACC;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hAACC;
defparam \readdata~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hAACC;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~10 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hAACC;
defparam \readdata~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hAACC;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hAACC;
defparam \readdata~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hAACC;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hAACC;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hAACC;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hAACC;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hAACC;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hAACC;
defparam \readdata~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~20 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hAACC;
defparam \readdata~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~21 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hAACC;
defparam \readdata~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~23 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~23_combout ),
	.cout());
defparam \readdata~23 .lut_mask = 16'hAACC;
defparam \readdata~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~24 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~24_combout ),
	.cout());
defparam \readdata~24 .lut_mask = 16'hAACC;
defparam \readdata~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~25 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~25_combout ),
	.cout());
defparam \readdata~25 .lut_mask = 16'hAACC;
defparam \readdata~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~26 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~26_combout ),
	.cout());
defparam \readdata~26 .lut_mask = 16'hAACC;
defparam \readdata~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~27 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hAACC;
defparam \readdata~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~28 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hAACC;
defparam \readdata~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~29 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~29_combout ),
	.cout());
defparam \readdata~29 .lut_mask = 16'hAACC;
defparam \readdata~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~30 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hAACC;
defparam \readdata~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~31 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~31_combout ),
	.cout());
defparam \readdata~31 .lut_mask = 16'hAACC;
defparam \readdata~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~32 (
	.dataa(\readdata~0_combout ),
	.datab(\the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.datac(gnd),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~32_combout ),
	.cout());
defparam \readdata~32 .lut_mask = 16'hAACC;
defparam \readdata~32 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_cpu_cpu_debug_slave_wrapper (
	sr_0,
	MonDReg_0,
	MonDReg_2,
	MonDReg_3,
	MonDReg_4,
	MonDReg_27,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_10,
	MonDReg_8,
	MonDReg_18,
	MonDReg_29,
	ir_out_0,
	ir_out_1,
	jdo_22,
	jdo_35,
	take_action_ocimem_a,
	jdo_34,
	take_action_ocimem_a1,
	break_readreg_0,
	hbreak_enabled,
	break_readreg_1,
	MonDReg_1,
	jdo_0,
	jdo_37,
	jdo_36,
	take_no_action_break_a,
	jdo_3,
	take_action_ocimem_b,
	monitor_ready,
	jdo_17,
	jdo_21,
	jdo_20,
	break_readreg_21,
	MonDReg_21,
	monitor_error,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_19,
	jdo_18,
	break_readreg_22,
	MonDReg_22,
	jdo_24,
	break_readreg_3,
	jdo_2,
	jdo_5,
	break_readreg_16,
	MonDReg_16,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	jdo_23,
	break_readreg_23,
	MonDReg_23,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	break_readreg_26,
	MonDReg_26,
	break_readreg_24,
	MonDReg_24,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_9,
	MonDReg_7,
	MonDReg_6,
	MonDReg_17,
	MonDReg_28,
	MonDReg_31,
	MonDReg_30,
	break_readreg_17,
	jdo_16,
	resetlatch,
	break_readreg_31,
	break_readreg_30,
	break_readreg_29,
	break_readreg_28,
	break_readreg_18,
	jdo_7,
	break_readreg_5,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_6,
	break_readreg_15,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
input 	MonDReg_2;
input 	MonDReg_3;
input 	MonDReg_4;
input 	MonDReg_27;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_10;
input 	MonDReg_8;
input 	MonDReg_18;
input 	MonDReg_29;
output 	ir_out_0;
output 	ir_out_1;
output 	jdo_22;
output 	jdo_35;
output 	take_action_ocimem_a;
output 	jdo_34;
output 	take_action_ocimem_a1;
input 	break_readreg_0;
input 	hbreak_enabled;
input 	break_readreg_1;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_37;
output 	jdo_36;
output 	take_no_action_break_a;
output 	jdo_3;
output 	take_action_ocimem_b;
input 	monitor_ready;
output 	jdo_17;
output 	jdo_21;
output 	jdo_20;
input 	break_readreg_21;
input 	MonDReg_21;
input 	monitor_error;
input 	break_readreg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
output 	jdo_19;
output 	jdo_18;
input 	break_readreg_22;
input 	MonDReg_22;
output 	jdo_24;
input 	break_readreg_3;
output 	jdo_2;
output 	jdo_5;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	jdo_23;
input 	break_readreg_23;
input 	MonDReg_23;
input 	break_readreg_4;
output 	jdo_6;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_24;
input 	MonDReg_24;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_9;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_17;
input 	MonDReg_28;
input 	MonDReg_31;
input 	MonDReg_30;
input 	break_readreg_17;
output 	jdo_16;
input 	resetlatch;
input 	break_readreg_31;
input 	break_readreg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	break_readreg_18;
output 	jdo_7;
input 	break_readreg_5;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	break_readreg_6;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[35]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[31]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[7]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[15]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[1]~q ;
wire \usb_system_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \usb_system_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[2]~q ;
wire \usb_system_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[22]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[34]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[3]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[23]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[36]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[4]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[37]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[17]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[21]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[20]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[24]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[5]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[26]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[28]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[27]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[25]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[18]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[33]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[32]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[30]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[29]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[19]~q ;
wire \usb_system_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[6]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[16]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[8]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[14]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[13]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[12]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[11]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[10]~q ;
wire \the_usb_system_cpu_cpu_debug_slave_tck|sr[9]~q ;


usb_system_sld_virtual_jtag_basic_1 usb_system_cpu_cpu_debug_slave_phy(
	.virtual_state_cdr1(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.virtual_state_udr(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

usb_system_usb_system_cpu_cpu_debug_slave_sysclk the_usb_system_cpu_cpu_debug_slave_sysclk(
	.sr_0(sr_0),
	.sr_35(\the_usb_system_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_usb_system_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.sr_7(\the_usb_system_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_usb_system_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.sr_1(\the_usb_system_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.jdo_22(jdo_22),
	.jdo_35(jdo_35),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_34(jdo_34),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.sr_2(\the_usb_system_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.virtual_state_uir(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_22(\the_usb_system_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.sr_34(\the_usb_system_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_3(\the_usb_system_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.jdo_0(jdo_0),
	.jdo_37(jdo_37),
	.jdo_36(jdo_36),
	.take_no_action_break_a(take_no_action_break_a),
	.jdo_3(jdo_3),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.jdo_17(jdo_17),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.sr_23(\the_usb_system_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.sr_36(\the_usb_system_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_4(\the_usb_system_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_37(\the_usb_system_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_25(jdo_25),
	.sr_17(\the_usb_system_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.jdo_33(jdo_33),
	.jdo_32(jdo_32),
	.jdo_31(jdo_31),
	.jdo_30(jdo_30),
	.jdo_29(jdo_29),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.sr_21(\the_usb_system_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_usb_system_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_24(\the_usb_system_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.jdo_24(jdo_24),
	.sr_5(\the_usb_system_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.sr_26(\the_usb_system_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_usb_system_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_usb_system_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_usb_system_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.sr_18(\the_usb_system_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.sr_33(\the_usb_system_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_usb_system_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_usb_system_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_usb_system_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.sr_19(\the_usb_system_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.jdo_23(jdo_23),
	.virtual_state_udr(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.sr_6(\the_usb_system_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.jdo_6(jdo_6),
	.jdo_16(jdo_16),
	.jdo_7(jdo_7),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_8(jdo_8),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_11(jdo_11),
	.jdo_10(jdo_10),
	.jdo_9(jdo_9),
	.sr_16(\the_usb_system_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.sr_8(\the_usb_system_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.sr_14(\the_usb_system_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_usb_system_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_usb_system_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_usb_system_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_usb_system_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_usb_system_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

usb_system_usb_system_cpu_cpu_debug_slave_tck the_usb_system_cpu_cpu_debug_slave_tck(
	.sr_0(sr_0),
	.MonDReg_0(MonDReg_0),
	.sr_35(\the_usb_system_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.MonDReg_2(MonDReg_2),
	.MonDReg_3(MonDReg_3),
	.sr_31(\the_usb_system_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.MonDReg_4(MonDReg_4),
	.MonDReg_27(MonDReg_27),
	.MonDReg_11(MonDReg_11),
	.MonDReg_12(MonDReg_12),
	.MonDReg_5(MonDReg_5),
	.MonDReg_10(MonDReg_10),
	.MonDReg_8(MonDReg_8),
	.MonDReg_18(MonDReg_18),
	.MonDReg_29(MonDReg_29),
	.sr_7(\the_usb_system_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_usb_system_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.sr_1(\the_usb_system_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.virtual_state_cdr(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.sr_2(\the_usb_system_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.virtual_state_uir(\usb_system_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.hbreak_enabled(hbreak_enabled),
	.sr_22(\the_usb_system_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.sr_34(\the_usb_system_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_3(\the_usb_system_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.monitor_ready(monitor_ready),
	.sr_23(\the_usb_system_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.MonDReg_21(MonDReg_21),
	.sr_36(\the_usb_system_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.monitor_error(monitor_error),
	.sr_4(\the_usb_system_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.sr_37(\the_usb_system_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.sr_17(\the_usb_system_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.sr_21(\the_usb_system_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_usb_system_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_24(\the_usb_system_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.MonDReg_22(MonDReg_22),
	.sr_5(\the_usb_system_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_26(\the_usb_system_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_usb_system_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_usb_system_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_usb_system_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.sr_18(\the_usb_system_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.sr_33(\the_usb_system_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_usb_system_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_usb_system_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_usb_system_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.sr_19(\the_usb_system_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.break_readreg_23(break_readreg_23),
	.MonDReg_23(MonDReg_23),
	.sr_6(\the_usb_system_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_27(break_readreg_27),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.MonDReg_15(MonDReg_15),
	.MonDReg_9(MonDReg_9),
	.MonDReg_7(MonDReg_7),
	.MonDReg_6(MonDReg_6),
	.MonDReg_17(MonDReg_17),
	.MonDReg_28(MonDReg_28),
	.MonDReg_31(MonDReg_31),
	.MonDReg_30(MonDReg_30),
	.break_readreg_17(break_readreg_17),
	.resetlatch(resetlatch),
	.break_readreg_31(break_readreg_31),
	.break_readreg_30(break_readreg_30),
	.break_readreg_29(break_readreg_29),
	.break_readreg_28(break_readreg_28),
	.break_readreg_18(break_readreg_18),
	.break_readreg_5(break_readreg_5),
	.sr_16(\the_usb_system_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.break_readreg_6(break_readreg_6),
	.sr_8(\the_usb_system_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.sr_14(\the_usb_system_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_usb_system_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_usb_system_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_usb_system_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_usb_system_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_usb_system_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_15(break_readreg_15),
	.break_readreg_7(break_readreg_7),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_10(break_readreg_10),
	.break_readreg_9(break_readreg_9),
	.break_readreg_8(break_readreg_8),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module usb_system_sld_virtual_jtag_basic_1 (
	virtual_state_cdr1,
	virtual_state_sdr,
	virtual_state_uir,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_cdr1;
output 	virtual_state_sdr;
output 	virtual_state_uir;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb virtual_state_cdr(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_3),
	.datad(splitter_nodes_receive_1_3),
	.cin(gnd),
	.combout(virtual_state_cdr1),
	.cout());
defparam virtual_state_cdr.lut_mask = 16'hAFFF;
defparam virtual_state_cdr.sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_sdr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_sdr),
	.cout());
defparam \virtual_state_sdr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_sdr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_uir~0 (
	.dataa(virtual_ir_scan_reg),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(virtual_state_uir),
	.cout());
defparam \virtual_state_uir~0 .lut_mask = 16'hFEFE;
defparam \virtual_state_uir~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_udr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_udr),
	.cout());
defparam \virtual_state_udr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_udr~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_cpu_cpu_debug_slave_sysclk (
	sr_0,
	sr_35,
	sr_31,
	sr_7,
	sr_15,
	sr_1,
	jdo_22,
	jdo_35,
	take_action_ocimem_a1,
	jdo_34,
	take_action_ocimem_a2,
	sr_2,
	virtual_state_uir,
	sr_22,
	sr_34,
	sr_3,
	jdo_0,
	jdo_37,
	jdo_36,
	take_no_action_break_a,
	jdo_3,
	take_action_ocimem_b1,
	jdo_17,
	jdo_21,
	jdo_20,
	sr_23,
	sr_36,
	sr_4,
	jdo_1,
	jdo_4,
	sr_37,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	sr_17,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_19,
	jdo_18,
	sr_21,
	sr_20,
	sr_24,
	jdo_24,
	sr_5,
	jdo_2,
	jdo_5,
	sr_26,
	sr_28,
	sr_27,
	sr_25,
	sr_18,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_19,
	jdo_23,
	virtual_state_udr,
	sr_6,
	jdo_6,
	jdo_16,
	jdo_7,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	sr_16,
	sr_8,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_0;
input 	sr_35;
input 	sr_31;
input 	sr_7;
input 	sr_15;
input 	sr_1;
output 	jdo_22;
output 	jdo_35;
output 	take_action_ocimem_a1;
output 	jdo_34;
output 	take_action_ocimem_a2;
input 	sr_2;
input 	virtual_state_uir;
input 	sr_22;
input 	sr_34;
input 	sr_3;
output 	jdo_0;
output 	jdo_37;
output 	jdo_36;
output 	take_no_action_break_a;
output 	jdo_3;
output 	take_action_ocimem_b1;
output 	jdo_17;
output 	jdo_21;
output 	jdo_20;
input 	sr_23;
input 	sr_36;
input 	sr_4;
output 	jdo_1;
output 	jdo_4;
input 	sr_37;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
input 	sr_17;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
output 	jdo_19;
output 	jdo_18;
input 	sr_21;
input 	sr_20;
input 	sr_24;
output 	jdo_24;
input 	sr_5;
output 	jdo_2;
output 	jdo_5;
input 	sr_26;
input 	sr_28;
input 	sr_27;
input 	sr_25;
input 	sr_18;
input 	sr_33;
input 	sr_32;
input 	sr_30;
input 	sr_29;
input 	sr_19;
output 	jdo_23;
input 	virtual_state_udr;
input 	sr_6;
output 	jdo_6;
output 	jdo_16;
output 	jdo_7;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	sr_16;
input 	sr_8;
input 	sr_14;
input 	sr_13;
input 	sr_12;
input 	sr_11;
input 	sr_10;
input 	sr_9;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \enable_action_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;
wire \ir[1]~q ;
wire \ir[0]~q ;


usb_system_altera_std_synchronizer_2 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_1 the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cycloneive_lcell_comb \take_action_ocimem_a~0 (
	.dataa(\enable_action_strobe~q ),
	.datab(gnd),
	.datac(\ir[1]~q ),
	.datad(\ir[0]~q ),
	.cin(gnd),
	.combout(take_action_ocimem_a1),
	.cout());
defparam \take_action_ocimem_a~0 .lut_mask = 16'hAFFF;
defparam \take_action_ocimem_a~0 .sum_lutc_input = "datac";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_a(
	.dataa(jdo_35),
	.datab(gnd),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(take_action_ocimem_a2),
	.cout());
defparam take_action_ocimem_a.lut_mask = 16'hFFF5;
defparam take_action_ocimem_a.sum_lutc_input = "datac";

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

cycloneive_lcell_comb \take_no_action_break_a~0 (
	.dataa(\ir[1]~q ),
	.datab(\enable_action_strobe~q ),
	.datac(gnd),
	.datad(\ir[0]~q ),
	.cin(gnd),
	.combout(take_no_action_break_a),
	.cout());
defparam \take_no_action_break_a~0 .lut_mask = 16'hEEFF;
defparam \take_no_action_break_a~0 .sum_lutc_input = "datac";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_b(
	.dataa(jdo_35),
	.datab(\enable_action_strobe~q ),
	.datac(\ir[1]~q ),
	.datad(\ir[0]~q ),
	.cin(gnd),
	.combout(take_action_ocimem_b1),
	.cout());
defparam take_action_ocimem_b.lut_mask = 16'hEFFF;
defparam take_action_ocimem_b.sum_lutc_input = "datac";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cycloneive_lcell_comb \update_jdo_strobe~0 (
	.dataa(\the_altera_std_synchronizer3|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_udr~q ),
	.cin(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.cout());
defparam \update_jdo_strobe~0 .lut_mask = 16'hAAFF;
defparam \update_jdo_strobe~0 .sum_lutc_input = "datac";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\enable_action_strobe~q ),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cycloneive_lcell_comb \jxuir~0 (
	.dataa(\the_altera_std_synchronizer4|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_uir~q ),
	.cin(gnd),
	.combout(\jxuir~0_combout ),
	.cout());
defparam \jxuir~0 .lut_mask = 16'hAAFF;
defparam \jxuir~0 .sum_lutc_input = "datac";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(\ir[1]~q ),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(\ir[0]~q ),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_1 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_2 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_usb_system_cpu_cpu_debug_slave_tck (
	sr_0,
	MonDReg_0,
	sr_35,
	MonDReg_2,
	MonDReg_3,
	sr_31,
	MonDReg_4,
	MonDReg_27,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_10,
	MonDReg_8,
	MonDReg_18,
	MonDReg_29,
	sr_7,
	sr_15,
	ir_out_0,
	ir_out_1,
	sr_1,
	virtual_state_cdr,
	virtual_state_sdr,
	sr_2,
	break_readreg_0,
	virtual_state_uir,
	hbreak_enabled,
	sr_22,
	sr_34,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	monitor_ready,
	sr_23,
	break_readreg_21,
	MonDReg_21,
	sr_36,
	monitor_error,
	sr_4,
	break_readreg_2,
	sr_37,
	sr_17,
	sr_21,
	sr_20,
	sr_24,
	break_readreg_22,
	MonDReg_22,
	sr_5,
	break_readreg_3,
	sr_26,
	sr_28,
	sr_27,
	sr_25,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_19,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	break_readreg_23,
	MonDReg_23,
	sr_6,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	break_readreg_26,
	MonDReg_26,
	break_readreg_24,
	MonDReg_24,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_9,
	MonDReg_7,
	MonDReg_6,
	MonDReg_17,
	MonDReg_28,
	MonDReg_31,
	MonDReg_30,
	break_readreg_17,
	resetlatch,
	break_readreg_31,
	break_readreg_30,
	break_readreg_29,
	break_readreg_28,
	break_readreg_18,
	break_readreg_5,
	sr_16,
	break_readreg_6,
	sr_8,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	break_readreg_15,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
output 	sr_35;
input 	MonDReg_2;
input 	MonDReg_3;
output 	sr_31;
input 	MonDReg_4;
input 	MonDReg_27;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_10;
input 	MonDReg_8;
input 	MonDReg_18;
input 	MonDReg_29;
output 	sr_7;
output 	sr_15;
output 	ir_out_0;
output 	ir_out_1;
output 	sr_1;
input 	virtual_state_cdr;
input 	virtual_state_sdr;
output 	sr_2;
input 	break_readreg_0;
input 	virtual_state_uir;
input 	hbreak_enabled;
output 	sr_22;
output 	sr_34;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
input 	monitor_ready;
output 	sr_23;
input 	break_readreg_21;
input 	MonDReg_21;
output 	sr_36;
input 	monitor_error;
output 	sr_4;
input 	break_readreg_2;
output 	sr_37;
output 	sr_17;
output 	sr_21;
output 	sr_20;
output 	sr_24;
input 	break_readreg_22;
input 	MonDReg_22;
output 	sr_5;
input 	break_readreg_3;
output 	sr_26;
output 	sr_28;
output 	sr_27;
output 	sr_25;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
output 	sr_33;
output 	sr_32;
output 	sr_30;
output 	sr_29;
output 	sr_19;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	break_readreg_23;
input 	MonDReg_23;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_24;
input 	MonDReg_24;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_9;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_17;
input 	MonDReg_28;
input 	MonDReg_31;
input 	MonDReg_30;
input 	break_readreg_17;
input 	resetlatch;
input 	break_readreg_31;
input 	break_readreg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	break_readreg_18;
input 	break_readreg_5;
output 	sr_16;
input 	break_readreg_6;
output 	sr_8;
output 	sr_14;
output 	sr_13;
output 	sr_12;
output 	sr_11;
output 	sr_10;
output 	sr_9;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \DRsize.000~q ;
wire \sr[0]~5_combout ;
wire \Mux37~0_combout ;
wire \sr~10_combout ;
wire \DRsize.100~q ;
wire \sr[35]~6_combout ;
wire \sr~20_combout ;
wire \sr~21_combout ;
wire \sr~22_combout ;
wire \sr[31]~56_combout ;
wire \sr[31]~7_combout ;
wire \Mux30~0_combout ;
wire \sr[7]~8_combout ;
wire \sr[29]~83_combout ;
wire \DRsize.010~q ;
wire \sr[15]~9_combout ;
wire \sr~71_combout ;
wire \sr~72_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr[2]~13_combout ;
wire \sr~14_combout ;
wire \sr~15_combout ;
wire \sr~16_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr[29]~19_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr[37]~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~50_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~55_combout ;
wire \sr~57_combout ;
wire \sr~58_combout ;
wire \sr~59_combout ;
wire \sr~60_combout ;
wire \sr~61_combout ;
wire \sr~62_combout ;
wire \sr~63_combout ;
wire \sr~64_combout ;
wire \sr~65_combout ;
wire \sr~66_combout ;
wire \sr~67_combout ;
wire \sr~68_combout ;
wire \sr~69_combout ;
wire \sr~70_combout ;
wire \sr~73_combout ;
wire \sr~74_combout ;
wire \sr~75_combout ;
wire \sr~76_combout ;
wire \sr~77_combout ;
wire \sr~78_combout ;
wire \sr~79_combout ;
wire \sr~80_combout ;
wire \sr~81_combout ;
wire \sr~82_combout ;


usb_system_altera_std_synchronizer_4 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

usb_system_altera_std_synchronizer_3 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr[0]~5_combout ),
	.asdata(\sr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr[35]~6_combout ),
	.asdata(\sr~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr[31]~7_combout ),
	.asdata(sr_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr[7]~8_combout ),
	.asdata(sr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr[15]~9_combout ),
	.asdata(\sr~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~29_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~29_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[2]~13_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cycloneive_lcell_comb \sr[0]~5 (
	.dataa(altera_internal_jtag1),
	.datab(sr_1),
	.datac(gnd),
	.datad(\DRsize.000~q ),
	.cin(gnd),
	.combout(\sr[0]~5_combout ),
	.cout());
defparam \sr[0]~5 .lut_mask = 16'hAACC;
defparam \sr[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux37~0 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
defparam \Mux37~0 .lut_mask = 16'h7777;
defparam \Mux37~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~10 (
	.dataa(sr_0),
	.datab(virtual_state_cdr),
	.datac(\the_altera_std_synchronizer2|dreg[0]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~10_combout ),
	.cout());
defparam \sr~10 .lut_mask = 16'hFFB8;
defparam \sr~10 .sum_lutc_input = "datac";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cycloneive_lcell_comb \sr[35]~6 (
	.dataa(sr_36),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.100~q ),
	.cin(gnd),
	.combout(\sr[35]~6_combout ),
	.cout());
defparam \sr[35]~6 .lut_mask = 16'hAACC;
defparam \sr[35]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~20 (
	.dataa(irf_reg_1_2),
	.datab(state_3),
	.datac(splitter_nodes_receive_1_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~20_combout ),
	.cout());
defparam \sr~20 .lut_mask = 16'hFDFF;
defparam \sr~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~21 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(sr_35),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr~21_combout ),
	.cout());
defparam \sr~21 .lut_mask = 16'hFFFE;
defparam \sr~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~22 (
	.dataa(irf_reg_0_2),
	.datab(\the_altera_std_synchronizer1|dreg[0]~q ),
	.datac(\sr~20_combout ),
	.datad(\sr~21_combout ),
	.cin(gnd),
	.combout(\sr~22_combout ),
	.cout());
defparam \sr~22 .lut_mask = 16'hFFFD;
defparam \sr~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~56 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(break_readreg_30),
	.datad(MonDReg_30),
	.cin(gnd),
	.combout(\sr[31]~56_combout ),
	.cout());
defparam \sr[31]~56 .lut_mask = 16'hFFF6;
defparam \sr[31]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~7 (
	.dataa(sr_31),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(\sr[31]~56_combout ),
	.cin(gnd),
	.combout(\sr[31]~7_combout ),
	.cout());
defparam \sr[31]~7 .lut_mask = 16'hBF8F;
defparam \sr[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~0 (
	.dataa(break_readreg_6),
	.datab(MonDReg_6),
	.datac(irf_reg_1_2),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hACFF;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[7]~8 (
	.dataa(\Mux30~0_combout ),
	.datab(sr_7),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr[7]~8_combout ),
	.cout());
defparam \sr[7]~8 .lut_mask = 16'hAACC;
defparam \sr[7]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[29]~83 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sr[29]~83_combout ),
	.cout());
defparam \sr[29]~83 .lut_mask = 16'hEEEE;
defparam \sr[29]~83 .sum_lutc_input = "datac";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[29]~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cycloneive_lcell_comb \sr[15]~9 (
	.dataa(sr_16),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.010~q ),
	.cin(gnd),
	.combout(\sr[15]~9_combout ),
	.cout());
defparam \sr[15]~9 .lut_mask = 16'hAACC;
defparam \sr[15]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~71 (
	.dataa(break_readreg_14),
	.datab(MonDReg_14),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~71_combout ),
	.cout());
defparam \sr~71 .lut_mask = 16'hAACC;
defparam \sr~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~72 (
	.dataa(sr_15),
	.datab(virtual_state_cdr),
	.datac(\sr~71_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~72_combout ),
	.cout());
defparam \sr~72 .lut_mask = 16'hB8FF;
defparam \sr~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~11 (
	.dataa(break_readreg_0),
	.datab(MonDReg_0),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~11_combout ),
	.cout());
defparam \sr~11 .lut_mask = 16'hAACC;
defparam \sr~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~12 (
	.dataa(sr_2),
	.datab(virtual_state_sdr),
	.datac(\sr~11_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~12_combout ),
	.cout());
defparam \sr~12 .lut_mask = 16'hB8FF;
defparam \sr~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[2]~13 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr[2]~13_combout ),
	.cout());
defparam \sr[2]~13 .lut_mask = 16'hFEFF;
defparam \sr[2]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~14 (
	.dataa(break_readreg_1),
	.datab(MonDReg_1),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~14_combout ),
	.cout());
defparam \sr~14 .lut_mask = 16'hAACC;
defparam \sr~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~15 (
	.dataa(sr_3),
	.datab(virtual_state_sdr),
	.datac(\sr~14_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~15_combout ),
	.cout());
defparam \sr~15 .lut_mask = 16'hB8FF;
defparam \sr~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~16 (
	.dataa(break_readreg_21),
	.datab(MonDReg_21),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~16_combout ),
	.cout());
defparam \sr~16 .lut_mask = 16'hAACC;
defparam \sr~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~17 (
	.dataa(virtual_state_sdr),
	.datab(irf_reg_0_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~17_combout ),
	.cout());
defparam \sr~17 .lut_mask = 16'hEEFF;
defparam \sr~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~18 (
	.dataa(virtual_state_sdr),
	.datab(sr_23),
	.datac(\sr~16_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~18_combout ),
	.cout());
defparam \sr~18 .lut_mask = 16'hFEFF;
defparam \sr~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[29]~19 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[29]~19_combout ),
	.cout());
defparam \sr[29]~19 .lut_mask = 16'hFF7F;
defparam \sr[29]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~23 (
	.dataa(sr_35),
	.datab(virtual_state_sdr),
	.datac(monitor_error),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~23_combout ),
	.cout());
defparam \sr~23 .lut_mask = 16'hFFB8;
defparam \sr~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~24 (
	.dataa(break_readreg_2),
	.datab(MonDReg_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~24_combout ),
	.cout());
defparam \sr~24 .lut_mask = 16'hAACC;
defparam \sr~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~25 (
	.dataa(sr_4),
	.datab(virtual_state_sdr),
	.datac(\sr~24_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~25_combout ),
	.cout());
defparam \sr~25 .lut_mask = 16'hB8FF;
defparam \sr~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~26 (
	.dataa(break_readreg_22),
	.datab(MonDReg_22),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~26_combout ),
	.cout());
defparam \sr~26 .lut_mask = 16'hAACC;
defparam \sr~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~27 (
	.dataa(virtual_state_sdr),
	.datab(sr_24),
	.datac(\sr~26_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~27_combout ),
	.cout());
defparam \sr~27 .lut_mask = 16'hFEFF;
defparam \sr~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~28 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(sr_37),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~28_combout ),
	.cout());
defparam \sr~28 .lut_mask = 16'hFEFF;
defparam \sr~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[37]~29 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[37]~29_combout ),
	.cout());
defparam \sr[37]~29 .lut_mask = 16'hFF7D;
defparam \sr[37]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~30 (
	.dataa(break_readreg_3),
	.datab(MonDReg_3),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~30_combout ),
	.cout());
defparam \sr~30 .lut_mask = 16'hAACC;
defparam \sr~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~31 (
	.dataa(sr_5),
	.datab(virtual_state_sdr),
	.datac(\sr~30_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~31_combout ),
	.cout());
defparam \sr~31 .lut_mask = 16'hB8FF;
defparam \sr~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~32 (
	.dataa(altera_internal_jtag1),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~32_combout ),
	.cout());
defparam \sr~32 .lut_mask = 16'hFEFF;
defparam \sr~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~33 (
	.dataa(break_readreg_16),
	.datab(MonDReg_16),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~33_combout ),
	.cout());
defparam \sr~33 .lut_mask = 16'hAACC;
defparam \sr~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~34 (
	.dataa(virtual_state_sdr),
	.datab(sr_18),
	.datac(\sr~33_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~34_combout ),
	.cout());
defparam \sr~34 .lut_mask = 16'hFEFF;
defparam \sr~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~35 (
	.dataa(break_readreg_20),
	.datab(MonDReg_20),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~35_combout ),
	.cout());
defparam \sr~35 .lut_mask = 16'hAACC;
defparam \sr~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~36 (
	.dataa(virtual_state_sdr),
	.datab(sr_22),
	.datac(\sr~35_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~36_combout ),
	.cout());
defparam \sr~36 .lut_mask = 16'hFEFF;
defparam \sr~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~37 (
	.dataa(break_readreg_19),
	.datab(MonDReg_19),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~37_combout ),
	.cout());
defparam \sr~37 .lut_mask = 16'hAACC;
defparam \sr~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~38 (
	.dataa(virtual_state_sdr),
	.datab(sr_21),
	.datac(\sr~37_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~38_combout ),
	.cout());
defparam \sr~38 .lut_mask = 16'hFEFF;
defparam \sr~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~39 (
	.dataa(break_readreg_23),
	.datab(MonDReg_23),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~39_combout ),
	.cout());
defparam \sr~39 .lut_mask = 16'hAACC;
defparam \sr~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~40 (
	.dataa(virtual_state_sdr),
	.datab(sr_25),
	.datac(\sr~39_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~40_combout ),
	.cout());
defparam \sr~40 .lut_mask = 16'hFEFF;
defparam \sr~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~41 (
	.dataa(break_readreg_4),
	.datab(MonDReg_4),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~41_combout ),
	.cout());
defparam \sr~41 .lut_mask = 16'hAACC;
defparam \sr~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~42 (
	.dataa(sr_6),
	.datab(virtual_state_sdr),
	.datac(\sr~41_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~42_combout ),
	.cout());
defparam \sr~42 .lut_mask = 16'hB8FF;
defparam \sr~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~43 (
	.dataa(break_readreg_25),
	.datab(MonDReg_25),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~43_combout ),
	.cout());
defparam \sr~43 .lut_mask = 16'hAACC;
defparam \sr~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~44 (
	.dataa(virtual_state_sdr),
	.datab(sr_27),
	.datac(\sr~43_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~44_combout ),
	.cout());
defparam \sr~44 .lut_mask = 16'hFEFF;
defparam \sr~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~45 (
	.dataa(break_readreg_27),
	.datab(MonDReg_27),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~45_combout ),
	.cout());
defparam \sr~45 .lut_mask = 16'hAACC;
defparam \sr~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~46 (
	.dataa(virtual_state_sdr),
	.datab(sr_29),
	.datac(\sr~45_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~46_combout ),
	.cout());
defparam \sr~46 .lut_mask = 16'hFEFF;
defparam \sr~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~47 (
	.dataa(break_readreg_26),
	.datab(MonDReg_26),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~47_combout ),
	.cout());
defparam \sr~47 .lut_mask = 16'hAACC;
defparam \sr~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~48 (
	.dataa(virtual_state_sdr),
	.datab(sr_28),
	.datac(\sr~47_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~48_combout ),
	.cout());
defparam \sr~48 .lut_mask = 16'hFEFF;
defparam \sr~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~49 (
	.dataa(break_readreg_24),
	.datab(MonDReg_24),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~49_combout ),
	.cout());
defparam \sr~49 .lut_mask = 16'hAACC;
defparam \sr~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~50 (
	.dataa(virtual_state_sdr),
	.datab(sr_26),
	.datac(\sr~49_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~50_combout ),
	.cout());
defparam \sr~50 .lut_mask = 16'hFEFF;
defparam \sr~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~51 (
	.dataa(break_readreg_17),
	.datab(MonDReg_17),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~51_combout ),
	.cout());
defparam \sr~51 .lut_mask = 16'hAACC;
defparam \sr~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~52 (
	.dataa(virtual_state_sdr),
	.datab(sr_19),
	.datac(\sr~51_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~52_combout ),
	.cout());
defparam \sr~52 .lut_mask = 16'hFEFF;
defparam \sr~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~53 (
	.dataa(sr_34),
	.datab(virtual_state_sdr),
	.datac(resetlatch),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~53_combout ),
	.cout());
defparam \sr~53 .lut_mask = 16'hFFB8;
defparam \sr~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~54 (
	.dataa(break_readreg_31),
	.datab(MonDReg_31),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~54_combout ),
	.cout());
defparam \sr~54 .lut_mask = 16'hAACC;
defparam \sr~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~55 (
	.dataa(virtual_state_sdr),
	.datab(sr_33),
	.datac(\sr~54_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~55_combout ),
	.cout());
defparam \sr~55 .lut_mask = 16'hFEFF;
defparam \sr~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~57 (
	.dataa(break_readreg_29),
	.datab(MonDReg_29),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~57_combout ),
	.cout());
defparam \sr~57 .lut_mask = 16'hAACC;
defparam \sr~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~58 (
	.dataa(virtual_state_sdr),
	.datab(sr_31),
	.datac(\sr~57_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~58_combout ),
	.cout());
defparam \sr~58 .lut_mask = 16'hFEFF;
defparam \sr~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~59 (
	.dataa(break_readreg_28),
	.datab(MonDReg_28),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~59_combout ),
	.cout());
defparam \sr~59 .lut_mask = 16'hAACC;
defparam \sr~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~60 (
	.dataa(virtual_state_sdr),
	.datab(sr_30),
	.datac(\sr~59_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~60_combout ),
	.cout());
defparam \sr~60 .lut_mask = 16'hFEFF;
defparam \sr~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~61 (
	.dataa(break_readreg_18),
	.datab(MonDReg_18),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~61_combout ),
	.cout());
defparam \sr~61 .lut_mask = 16'hAACC;
defparam \sr~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~62 (
	.dataa(virtual_state_sdr),
	.datab(sr_20),
	.datac(\sr~61_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~62_combout ),
	.cout());
defparam \sr~62 .lut_mask = 16'hFEFF;
defparam \sr~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~63 (
	.dataa(break_readreg_5),
	.datab(MonDReg_5),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~63_combout ),
	.cout());
defparam \sr~63 .lut_mask = 16'hAACC;
defparam \sr~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~64 (
	.dataa(sr_7),
	.datab(virtual_state_sdr),
	.datac(\sr~63_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~64_combout ),
	.cout());
defparam \sr~64 .lut_mask = 16'hB8FF;
defparam \sr~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~65 (
	.dataa(break_readreg_15),
	.datab(MonDReg_15),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~65_combout ),
	.cout());
defparam \sr~65 .lut_mask = 16'hAACC;
defparam \sr~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~66 (
	.dataa(virtual_state_sdr),
	.datab(sr_17),
	.datac(\sr~65_combout ),
	.datad(\sr~17_combout ),
	.cin(gnd),
	.combout(\sr~66_combout ),
	.cout());
defparam \sr~66 .lut_mask = 16'hFEFF;
defparam \sr~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~67 (
	.dataa(break_readreg_7),
	.datab(MonDReg_7),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~67_combout ),
	.cout());
defparam \sr~67 .lut_mask = 16'hAACC;
defparam \sr~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~68 (
	.dataa(sr_9),
	.datab(virtual_state_sdr),
	.datac(\sr~67_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~68_combout ),
	.cout());
defparam \sr~68 .lut_mask = 16'hB8FF;
defparam \sr~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~69 (
	.dataa(break_readreg_13),
	.datab(MonDReg_13),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~69_combout ),
	.cout());
defparam \sr~69 .lut_mask = 16'hAACC;
defparam \sr~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~70 (
	.dataa(sr_15),
	.datab(virtual_state_sdr),
	.datac(\sr~69_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~70_combout ),
	.cout());
defparam \sr~70 .lut_mask = 16'hB8FF;
defparam \sr~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~73 (
	.dataa(break_readreg_12),
	.datab(MonDReg_12),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~73_combout ),
	.cout());
defparam \sr~73 .lut_mask = 16'hAACC;
defparam \sr~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~74 (
	.dataa(sr_14),
	.datab(virtual_state_sdr),
	.datac(\sr~73_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~74_combout ),
	.cout());
defparam \sr~74 .lut_mask = 16'hB8FF;
defparam \sr~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~75 (
	.dataa(break_readreg_11),
	.datab(MonDReg_11),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~75_combout ),
	.cout());
defparam \sr~75 .lut_mask = 16'hAACC;
defparam \sr~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~76 (
	.dataa(sr_13),
	.datab(virtual_state_sdr),
	.datac(\sr~75_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~76_combout ),
	.cout());
defparam \sr~76 .lut_mask = 16'hB8FF;
defparam \sr~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~77 (
	.dataa(break_readreg_10),
	.datab(MonDReg_10),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~77_combout ),
	.cout());
defparam \sr~77 .lut_mask = 16'hAACC;
defparam \sr~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~78 (
	.dataa(sr_12),
	.datab(virtual_state_sdr),
	.datac(\sr~77_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~78_combout ),
	.cout());
defparam \sr~78 .lut_mask = 16'hB8FF;
defparam \sr~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~79 (
	.dataa(break_readreg_9),
	.datab(MonDReg_9),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~79_combout ),
	.cout());
defparam \sr~79 .lut_mask = 16'hAACC;
defparam \sr~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~80 (
	.dataa(sr_11),
	.datab(virtual_state_sdr),
	.datac(\sr~79_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~80_combout ),
	.cout());
defparam \sr~80 .lut_mask = 16'hB8FF;
defparam \sr~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~81 (
	.dataa(break_readreg_8),
	.datab(MonDReg_8),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~81_combout ),
	.cout());
defparam \sr~81 .lut_mask = 16'hAACC;
defparam \sr~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~82 (
	.dataa(sr_10),
	.datab(virtual_state_sdr),
	.datac(\sr~81_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~82_combout ),
	.cout());
defparam \sr~82 .lut_mask = 16'hB8FF;
defparam \sr~82 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_4 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_usb_system_cpu_cpu_nios2_avalon_reg (
	r_sync_rst,
	address_8,
	oci_ienable_6,
	oci_ienable_5,
	oci_single_step_mode1,
	ociram_wr_en,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	Equal0,
	Equal01,
	take_action_ocireg,
	writedata_6,
	writedata_5,
	writedata_3,
	oci_ienable_22,
	Equal02,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	address_8;
output 	oci_ienable_6;
output 	oci_ienable_5;
output 	oci_single_step_mode1;
input 	ociram_wr_en;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
output 	Equal0;
output 	Equal01;
output 	take_action_ocireg;
input 	writedata_6;
input 	writedata_5;
input 	writedata_3;
output 	oci_ienable_22;
output 	Equal02;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \oci_ienable[6]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[5]~1_combout ;
wire \oci_single_step_mode~0_combout ;


dffeas \oci_ienable[6] (
	.clk(clk_clk),
	.d(\oci_ienable[6]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_6),
	.prn(vcc));
defparam \oci_ienable[6] .is_wysiwyg = "true";
defparam \oci_ienable[6] .power_up = "low";

dffeas \oci_ienable[5] (
	.clk(clk_clk),
	.d(\oci_ienable[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_5),
	.prn(vcc));
defparam \oci_ienable[5] .is_wysiwyg = "true";
defparam \oci_ienable[5] .power_up = "low";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(address_8),
	.datab(address_5),
	.datac(address_6),
	.datad(address_7),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hBFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(address_1),
	.datab(address_2),
	.datac(address_3),
	.datad(address_4),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocireg~0 (
	.dataa(ociram_wr_en),
	.datab(Equal0),
	.datac(Equal01),
	.datad(address_0),
	.cin(gnd),
	.combout(take_action_ocireg),
	.cout());
defparam \take_action_ocireg~0 .lut_mask = 16'hFEFF;
defparam \take_action_ocireg~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[22] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_22),
	.prn(vcc));
defparam \oci_ienable[22] .is_wysiwyg = "true";
defparam \oci_ienable[22] .power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(Equal0),
	.datab(Equal01),
	.datac(gnd),
	.datad(address_0),
	.cin(gnd),
	.combout(Equal02),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[6]~0 (
	.dataa(writedata_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[6]~0_combout ),
	.cout());
defparam \oci_ienable[6]~0 .lut_mask = 16'h5555;
defparam \oci_ienable[6]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(ociram_wr_en),
	.datab(address_0),
	.datac(Equal0),
	.datad(Equal01),
	.cin(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.cout());
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 16'hFFFE;
defparam \take_action_oci_intr_mask_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[5]~1 (
	.dataa(writedata_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[5]~1_combout ),
	.cout());
defparam \oci_ienable[5]~1 .lut_mask = 16'h5555;
defparam \oci_ienable[5]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_single_step_mode~0 (
	.dataa(writedata_3),
	.datab(oci_single_step_mode1),
	.datac(gnd),
	.datad(take_action_ocireg),
	.cin(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.cout());
defparam \oci_single_step_mode~0 .lut_mask = 16'hAACC;
defparam \oci_single_step_mode~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_cpu_cpu_nios2_oci_break (
	jdo_22,
	break_readreg_0,
	break_readreg_1,
	jdo_0,
	jdo_37,
	jdo_36,
	take_no_action_break_a,
	jdo_3,
	jdo_17,
	jdo_21,
	jdo_20,
	break_readreg_21,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_19,
	jdo_18,
	break_readreg_22,
	jdo_24,
	break_readreg_3,
	jdo_2,
	jdo_5,
	break_readreg_16,
	break_readreg_20,
	break_readreg_19,
	jdo_23,
	break_readreg_23,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	break_readreg_27,
	break_readreg_26,
	break_readreg_24,
	break_readreg_17,
	jdo_16,
	break_readreg_31,
	break_readreg_30,
	break_readreg_29,
	break_readreg_28,
	break_readreg_18,
	jdo_7,
	break_readreg_5,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_6,
	break_readreg_15,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	jdo_22;
output 	break_readreg_0;
output 	break_readreg_1;
input 	jdo_0;
input 	jdo_37;
input 	jdo_36;
input 	take_no_action_break_a;
input 	jdo_3;
input 	jdo_17;
input 	jdo_21;
input 	jdo_20;
output 	break_readreg_21;
output 	break_readreg_2;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_25;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
input 	jdo_19;
input 	jdo_18;
output 	break_readreg_22;
input 	jdo_24;
output 	break_readreg_3;
input 	jdo_2;
input 	jdo_5;
output 	break_readreg_16;
output 	break_readreg_20;
output 	break_readreg_19;
input 	jdo_23;
output 	break_readreg_23;
output 	break_readreg_4;
input 	jdo_6;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_24;
output 	break_readreg_17;
input 	jdo_16;
output 	break_readreg_31;
output 	break_readreg_30;
output 	break_readreg_29;
output 	break_readreg_28;
output 	break_readreg_18;
input 	jdo_7;
output 	break_readreg_5;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
output 	break_readreg_6;
output 	break_readreg_15;
output 	break_readreg_7;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_10;
output 	break_readreg_9;
output 	break_readreg_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg~0_combout ;
wire \break_readreg~1_combout ;
wire \break_readreg~2_combout ;
wire \break_readreg~3_combout ;
wire \break_readreg~4_combout ;
wire \break_readreg~5_combout ;
wire \break_readreg~6_combout ;
wire \break_readreg~7_combout ;
wire \break_readreg~8_combout ;
wire \break_readreg~9_combout ;
wire \break_readreg~10_combout ;
wire \break_readreg~11_combout ;
wire \break_readreg~12_combout ;
wire \break_readreg~13_combout ;
wire \break_readreg~14_combout ;
wire \break_readreg~15_combout ;
wire \break_readreg~16_combout ;
wire \break_readreg~17_combout ;
wire \break_readreg~18_combout ;
wire \break_readreg~19_combout ;
wire \break_readreg~20_combout ;
wire \break_readreg~21_combout ;
wire \break_readreg~22_combout ;
wire \break_readreg~23_combout ;
wire \break_readreg~24_combout ;
wire \break_readreg~25_combout ;
wire \break_readreg~26_combout ;
wire \break_readreg~27_combout ;
wire \break_readreg~28_combout ;
wire \break_readreg~29_combout ;
wire \break_readreg~30_combout ;
wire \break_readreg~31_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(\break_readreg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(\break_readreg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(\break_readreg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(\break_readreg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(\break_readreg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(\break_readreg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(\break_readreg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(\break_readreg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(\break_readreg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(\break_readreg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(\break_readreg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(\break_readreg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(\break_readreg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(\break_readreg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(\break_readreg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(\break_readreg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(\break_readreg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(\break_readreg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(\break_readreg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(\break_readreg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(\break_readreg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(\break_readreg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(\break_readreg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(\break_readreg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(\break_readreg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(\break_readreg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(\break_readreg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(\break_readreg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(\break_readreg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(\break_readreg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(\break_readreg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(\break_readreg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

cycloneive_lcell_comb \break_readreg~0 (
	.dataa(jdo_0),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~0_combout ),
	.cout());
defparam \break_readreg~0 .lut_mask = 16'hFEFF;
defparam \break_readreg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~1 (
	.dataa(jdo_1),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~1_combout ),
	.cout());
defparam \break_readreg~1 .lut_mask = 16'hFEFF;
defparam \break_readreg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~2 (
	.dataa(jdo_21),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~2_combout ),
	.cout());
defparam \break_readreg~2 .lut_mask = 16'hFEFF;
defparam \break_readreg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~3 (
	.dataa(jdo_2),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~3_combout ),
	.cout());
defparam \break_readreg~3 .lut_mask = 16'hFEFF;
defparam \break_readreg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~4 (
	.dataa(jdo_22),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~4_combout ),
	.cout());
defparam \break_readreg~4 .lut_mask = 16'hFEFF;
defparam \break_readreg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~5 (
	.dataa(jdo_3),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~5_combout ),
	.cout());
defparam \break_readreg~5 .lut_mask = 16'hFEFF;
defparam \break_readreg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~6 (
	.dataa(jdo_16),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~6_combout ),
	.cout());
defparam \break_readreg~6 .lut_mask = 16'hFEFF;
defparam \break_readreg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~7 (
	.dataa(jdo_20),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~7_combout ),
	.cout());
defparam \break_readreg~7 .lut_mask = 16'hFEFF;
defparam \break_readreg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~8 (
	.dataa(jdo_19),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~8_combout ),
	.cout());
defparam \break_readreg~8 .lut_mask = 16'hFEFF;
defparam \break_readreg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~9 (
	.dataa(jdo_23),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~9_combout ),
	.cout());
defparam \break_readreg~9 .lut_mask = 16'hFEFF;
defparam \break_readreg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~10 (
	.dataa(jdo_4),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~10_combout ),
	.cout());
defparam \break_readreg~10 .lut_mask = 16'hFEFF;
defparam \break_readreg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~11 (
	.dataa(jdo_25),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~11_combout ),
	.cout());
defparam \break_readreg~11 .lut_mask = 16'hFEFF;
defparam \break_readreg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~12 (
	.dataa(jdo_27),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~12_combout ),
	.cout());
defparam \break_readreg~12 .lut_mask = 16'hFEFF;
defparam \break_readreg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~13 (
	.dataa(jdo_26),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~13_combout ),
	.cout());
defparam \break_readreg~13 .lut_mask = 16'hFEFF;
defparam \break_readreg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~14 (
	.dataa(jdo_24),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~14_combout ),
	.cout());
defparam \break_readreg~14 .lut_mask = 16'hFEFF;
defparam \break_readreg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~15 (
	.dataa(jdo_17),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~15_combout ),
	.cout());
defparam \break_readreg~15 .lut_mask = 16'hFEFF;
defparam \break_readreg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~16 (
	.dataa(jdo_31),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~16_combout ),
	.cout());
defparam \break_readreg~16 .lut_mask = 16'hFEFF;
defparam \break_readreg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~17 (
	.dataa(jdo_30),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~17_combout ),
	.cout());
defparam \break_readreg~17 .lut_mask = 16'hFEFF;
defparam \break_readreg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~18 (
	.dataa(jdo_29),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~18_combout ),
	.cout());
defparam \break_readreg~18 .lut_mask = 16'hFEFF;
defparam \break_readreg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~19 (
	.dataa(jdo_28),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~19_combout ),
	.cout());
defparam \break_readreg~19 .lut_mask = 16'hFEFF;
defparam \break_readreg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~20 (
	.dataa(jdo_18),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~20_combout ),
	.cout());
defparam \break_readreg~20 .lut_mask = 16'hFEFF;
defparam \break_readreg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~21 (
	.dataa(jdo_5),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~21_combout ),
	.cout());
defparam \break_readreg~21 .lut_mask = 16'hFEFF;
defparam \break_readreg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~22 (
	.dataa(jdo_6),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~22_combout ),
	.cout());
defparam \break_readreg~22 .lut_mask = 16'hFEFF;
defparam \break_readreg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~23 (
	.dataa(jdo_15),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~23_combout ),
	.cout());
defparam \break_readreg~23 .lut_mask = 16'hFEFF;
defparam \break_readreg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~24 (
	.dataa(jdo_7),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~24_combout ),
	.cout());
defparam \break_readreg~24 .lut_mask = 16'hFEFF;
defparam \break_readreg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~25 (
	.dataa(jdo_13),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~25_combout ),
	.cout());
defparam \break_readreg~25 .lut_mask = 16'hFEFF;
defparam \break_readreg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~26 (
	.dataa(jdo_14),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~26_combout ),
	.cout());
defparam \break_readreg~26 .lut_mask = 16'hFEFF;
defparam \break_readreg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~27 (
	.dataa(jdo_12),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~27_combout ),
	.cout());
defparam \break_readreg~27 .lut_mask = 16'hFEFF;
defparam \break_readreg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~28 (
	.dataa(jdo_11),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~28_combout ),
	.cout());
defparam \break_readreg~28 .lut_mask = 16'hFEFF;
defparam \break_readreg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~29 (
	.dataa(jdo_10),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~29_combout ),
	.cout());
defparam \break_readreg~29 .lut_mask = 16'hFEFF;
defparam \break_readreg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~30 (
	.dataa(jdo_9),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~30_combout ),
	.cout());
defparam \break_readreg~30 .lut_mask = 16'hFEFF;
defparam \break_readreg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~31 (
	.dataa(jdo_8),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~31_combout ),
	.cout());
defparam \break_readreg~31 .lut_mask = 16'hFEFF;
defparam \break_readreg~31 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_cpu_cpu_nios2_oci_debug (
	jtag_break1,
	r_sync_rst,
	resetrequest1,
	jdo_22,
	jdo_35,
	take_action_ocimem_a,
	jdo_34,
	take_action_ocimem_a1,
	monitor_ready1,
	jdo_21,
	jdo_20,
	monitor_error1,
	writedata_0,
	take_action_ocireg,
	jdo_25,
	jdo_19,
	jdo_18,
	monitor_go1,
	jdo_24,
	writedata_1,
	jdo_23,
	resetlatch1,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	jtag_break1;
input 	r_sync_rst;
output 	resetrequest1;
input 	jdo_22;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	take_action_ocimem_a1;
output 	monitor_ready1;
input 	jdo_21;
input 	jdo_20;
output 	monitor_error1;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_25;
input 	jdo_19;
input 	jdo_18;
output 	monitor_go1;
input 	jdo_24;
input 	writedata_1;
input 	jdo_23;
output 	resetlatch1;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \jtag_break~1_combout ;
wire \always1~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


usb_system_altera_std_synchronizer_5 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(\jtag_break~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas resetrequest(
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(resetrequest1),
	.prn(vcc));
defparam resetrequest.is_wysiwyg = "true";
defparam resetrequest.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cycloneive_lcell_comb \break_on_reset~0 (
	.dataa(jdo_19),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(jdo_18),
	.cin(gnd),
	.combout(\break_on_reset~0_combout ),
	.cout());
defparam \break_on_reset~0 .lut_mask = 16'hEEFF;
defparam \break_on_reset~0 .sum_lutc_input = "datac";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cycloneive_lcell_comb \jtag_break~0 (
	.dataa(jtag_break1),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(\the_altera_std_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\jtag_break~0_combout ),
	.cout());
defparam \jtag_break~0 .lut_mask = 16'hAACC;
defparam \jtag_break~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_break~1 (
	.dataa(jdo_21),
	.datab(jtag_break1),
	.datac(gnd),
	.datad(jdo_20),
	.cin(gnd),
	.combout(\jtag_break~1_combout ),
	.cout());
defparam \jtag_break~1 .lut_mask = 16'hEEFF;
defparam \jtag_break~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(take_action_ocimem_a),
	.datab(jdo_34),
	.datac(jdo_25),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_ready~0 (
	.dataa(monitor_ready1),
	.datab(writedata_0),
	.datac(take_action_ocireg),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_ready~0_combout ),
	.cout());
defparam \monitor_ready~0 .lut_mask = 16'hFEFF;
defparam \monitor_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_error~0 (
	.dataa(monitor_error1),
	.datab(take_action_ocireg),
	.datac(writedata_1),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_error~0_combout ),
	.cout());
defparam \monitor_error~0 .lut_mask = 16'hFEFF;
defparam \monitor_error~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_go~0 (
	.dataa(jdo_23),
	.datab(monitor_go1),
	.datac(take_action_ocimem_a1),
	.datad(state_1),
	.cin(gnd),
	.combout(\monitor_go~0_combout ),
	.cout());
defparam \monitor_go~0 .lut_mask = 16'hFEFF;
defparam \monitor_go~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \resetlatch~0 (
	.dataa(take_action_ocimem_a1),
	.datab(resetlatch1),
	.datac(\the_altera_std_synchronizer|dreg[0]~q ),
	.datad(jdo_24),
	.cin(gnd),
	.combout(\resetlatch~0_combout ),
	.cout());
defparam \resetlatch~0 .lut_mask = 16'hFDFF;
defparam \resetlatch~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_std_synchronizer_5 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_usb_system_cpu_cpu_nios2_ocimem (
	MonDReg_0,
	q_a_0,
	MonDReg_2,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_21,
	MonDReg_3,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_18,
	q_a_19,
	q_a_17,
	q_a_27,
	q_a_28,
	q_a_31,
	q_a_30,
	q_a_29,
	MonDReg_4,
	MonDReg_27,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_10,
	MonDReg_8,
	MonDReg_18,
	MonDReg_29,
	waitrequest1,
	jdo_22,
	jdo_35,
	take_action_ocimem_a,
	jdo_34,
	take_action_ocimem_a1,
	write,
	address_8,
	read,
	MonDReg_1,
	jdo_3,
	take_action_ocimem_b,
	jdo_17,
	jdo_21,
	jdo_20,
	MonDReg_21,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	debugaccess,
	ociram_wr_en,
	r_early_rst,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	byteenable_0,
	jdo_25,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	writedata_6,
	writedata_5,
	jdo_19,
	jdo_18,
	writedata_3,
	MonDReg_22,
	jdo_24,
	writedata_1,
	jdo_5,
	MonDReg_16,
	MonDReg_20,
	MonDReg_19,
	jdo_23,
	writedata_2,
	writedata_4,
	MonDReg_23,
	writedata_21,
	byteenable_2,
	jdo_6,
	MonDReg_25,
	MonDReg_26,
	MonDReg_24,
	writedata_22,
	writedata_23,
	writedata_24,
	byteenable_3,
	writedata_25,
	writedata_26,
	writedata_11,
	byteenable_1,
	MonDReg_13,
	writedata_13,
	writedata_16,
	writedata_12,
	MonDReg_14,
	writedata_14,
	MonDReg_15,
	writedata_15,
	writedata_10,
	MonDReg_9,
	writedata_9,
	writedata_8,
	MonDReg_7,
	writedata_7,
	MonDReg_6,
	writedata_20,
	writedata_18,
	writedata_19,
	MonDReg_17,
	writedata_17,
	writedata_27,
	MonDReg_28,
	writedata_28,
	MonDReg_31,
	writedata_31,
	MonDReg_30,
	writedata_30,
	writedata_29,
	jdo_16,
	jdo_7,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_0;
output 	q_a_0;
output 	MonDReg_2;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_21;
output 	MonDReg_3;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_18;
output 	q_a_19;
output 	q_a_17;
output 	q_a_27;
output 	q_a_28;
output 	q_a_31;
output 	q_a_30;
output 	q_a_29;
output 	MonDReg_4;
output 	MonDReg_27;
output 	MonDReg_11;
output 	MonDReg_12;
output 	MonDReg_5;
output 	MonDReg_10;
output 	MonDReg_8;
output 	MonDReg_18;
output 	MonDReg_29;
output 	waitrequest1;
input 	jdo_22;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	take_action_ocimem_a1;
input 	write;
input 	address_8;
input 	read;
output 	MonDReg_1;
input 	jdo_3;
input 	take_action_ocimem_b;
input 	jdo_17;
input 	jdo_21;
input 	jdo_20;
output 	MonDReg_21;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	debugaccess;
output 	ociram_wr_en;
input 	r_early_rst;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
input 	byteenable_0;
input 	jdo_25;
input 	jdo_33;
input 	jdo_32;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
input 	writedata_6;
input 	writedata_5;
input 	jdo_19;
input 	jdo_18;
input 	writedata_3;
output 	MonDReg_22;
input 	jdo_24;
input 	writedata_1;
input 	jdo_5;
output 	MonDReg_16;
output 	MonDReg_20;
output 	MonDReg_19;
input 	jdo_23;
input 	writedata_2;
input 	writedata_4;
output 	MonDReg_23;
input 	writedata_21;
input 	byteenable_2;
input 	jdo_6;
output 	MonDReg_25;
output 	MonDReg_26;
output 	MonDReg_24;
input 	writedata_22;
input 	writedata_23;
input 	writedata_24;
input 	byteenable_3;
input 	writedata_25;
input 	writedata_26;
input 	writedata_11;
input 	byteenable_1;
output 	MonDReg_13;
input 	writedata_13;
input 	writedata_16;
input 	writedata_12;
output 	MonDReg_14;
input 	writedata_14;
output 	MonDReg_15;
input 	writedata_15;
input 	writedata_10;
output 	MonDReg_9;
input 	writedata_9;
input 	writedata_8;
output 	MonDReg_7;
input 	writedata_7;
output 	MonDReg_6;
input 	writedata_20;
input 	writedata_18;
input 	writedata_19;
output 	MonDReg_17;
input 	writedata_17;
input 	writedata_27;
output 	MonDReg_28;
input 	writedata_28;
output 	MonDReg_31;
input 	writedata_31;
output 	MonDReg_30;
input 	writedata_30;
input 	writedata_29;
input 	jdo_16;
input 	jdo_7;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~1_combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[3]~3_combout ;
wire \ociram_wr_data[4]~4_combout ;
wire \ociram_wr_data[21]~5_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[22]~6_combout ;
wire \ociram_wr_data[23]~7_combout ;
wire \ociram_wr_data[24]~8_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[25]~9_combout ;
wire \ociram_wr_data[26]~10_combout ;
wire \ociram_wr_data[11]~11_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[13]~12_combout ;
wire \ociram_wr_data[16]~13_combout ;
wire \ociram_wr_data[12]~14_combout ;
wire \ociram_wr_data[5]~15_combout ;
wire \ociram_wr_data[14]~16_combout ;
wire \ociram_wr_data[15]~17_combout ;
wire \ociram_wr_data[10]~18_combout ;
wire \ociram_wr_data[9]~19_combout ;
wire \ociram_wr_data[8]~20_combout ;
wire \ociram_wr_data[7]~21_combout ;
wire \ociram_wr_data[6]~22_combout ;
wire \ociram_wr_data[20]~23_combout ;
wire \ociram_wr_data[18]~24_combout ;
wire \ociram_wr_data[19]~25_combout ;
wire \ociram_wr_data[17]~26_combout ;
wire \ociram_wr_data[27]~27_combout ;
wire \ociram_wr_data[28]~28_combout ;
wire \ociram_wr_data[31]~29_combout ;
wire \ociram_wr_data[30]~30_combout ;
wire \ociram_wr_data[29]~31_combout ;
wire \MonARegAddrInc[0]~0_combout ;
wire \MonAReg~0_combout ;
wire \MonAReg[2]~q ;
wire \MonARegAddrInc[0]~1 ;
wire \MonARegAddrInc[1]~2_combout ;
wire \MonAReg~2_combout ;
wire \MonAReg[3]~q ;
wire \MonARegAddrInc[1]~3 ;
wire \MonARegAddrInc[2]~4_combout ;
wire \MonAReg~1_combout ;
wire \MonAReg[4]~q ;
wire \Equal0~0_combout ;
wire \MonAReg~3_combout ;
wire \MonAReg[10]~q ;
wire \MonARegAddrInc[2]~5 ;
wire \MonARegAddrInc[3]~6_combout ;
wire \MonAReg~8_combout ;
wire \MonAReg[5]~q ;
wire \MonARegAddrInc[3]~7 ;
wire \MonARegAddrInc[4]~8_combout ;
wire \MonAReg~7_combout ;
wire \MonAReg[6]~q ;
wire \MonARegAddrInc[4]~9 ;
wire \MonARegAddrInc[5]~10_combout ;
wire \MonAReg~6_combout ;
wire \MonAReg[7]~q ;
wire \MonARegAddrInc[5]~11 ;
wire \MonARegAddrInc[6]~12_combout ;
wire \MonAReg~5_combout ;
wire \MonAReg[8]~q ;
wire \MonARegAddrInc[6]~13 ;
wire \MonARegAddrInc[7]~14_combout ;
wire \MonAReg~4_combout ;
wire \MonAReg[9]~q ;
wire \MonARegAddrInc[7]~15 ;
wire \MonARegAddrInc[8]~16_combout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~1_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[0]~0_combout ;
wire \jtag_rd~0_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~12_combout ;
wire \MonDReg[2]~1_combout ;
wire \MonDReg[3]~2_combout ;
wire \MonDReg[4]~3_combout ;
wire \cfgrom_readdata[27]~0_combout ;
wire \MonDReg[27]~4_combout ;
wire \MonDReg[27]~21_combout ;
wire \MonDReg[11]~6_combout ;
wire \MonDReg[12]~7_combout ;
wire \Equal0~1_combout ;
wire \MonDReg[5]~5_combout ;
wire \MonDReg[10]~11_combout ;
wire \cfgrom_readdata[8]~1_combout ;
wire \MonDReg[8]~10_combout ;
wire \Equal0~2_combout ;
wire \MonDReg[18]~8_combout ;
wire \Equal0~3_combout ;
wire \MonDReg[29]~9_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~1_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~1_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~20_combout ;
wire \MonDReg~22_combout ;
wire \MonDReg~23_combout ;
wire \MonDReg~24_combout ;
wire \MonDReg~25_combout ;
wire \MonDReg~26_combout ;
wire \MonDReg~27_combout ;
wire \MonDReg~28_combout ;
wire \MonDReg~29_combout ;
wire \MonDReg~30_combout ;
wire \MonDReg~31_combout ;
wire \MonDReg~32_combout ;
wire \MonDReg~33_combout ;


usb_system_usb_system_cpu_cpu_ociram_sp_ram_module usb_system_cpu_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_21(q_a_21),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_20(q_a_20),
	.q_a_18(q_a_18),
	.q_a_19(q_a_19),
	.q_a_17(q_a_17),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_31(q_a_31),
	.q_a_30(q_a_30),
	.q_a_29(q_a_29),
	.ociram_wr_en(\ociram_wr_en~1_combout ),
	.r_early_rst(r_early_rst),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~3_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~4_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~5_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~6_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~7_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~8_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~9_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~10_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~11_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~12_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~13_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~14_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~15_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~16_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~17_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~18_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~19_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~20_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~21_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~22_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~23_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~24_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~25_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~26_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~27_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~28_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~29_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~30_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cycloneive_lcell_comb \ociram_wr_en~1 (
	.dataa(\jtag_ram_wr~q ),
	.datab(\jtag_ram_access~q ),
	.datac(ociram_wr_en),
	.datad(address_8),
	.cin(gnd),
	.combout(\ociram_wr_en~1_combout ),
	.cout());
defparam \ociram_wr_en~1 .lut_mask = 16'hB8FF;
defparam \ociram_wr_en~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(MonDReg_0),
	.datab(writedata_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.cout());
defparam \ociram_wr_data[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(address_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.cout());
defparam \ociram_addr[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_addr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[1]~1 (
	.dataa(\MonAReg[3]~q ),
	.datab(address_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.cout());
defparam \ociram_addr[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_addr[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[2]~2 (
	.dataa(\MonAReg[4]~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.cout());
defparam \ociram_addr[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_addr[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[3]~3 (
	.dataa(\MonAReg[5]~q ),
	.datab(address_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.cout());
defparam \ociram_addr[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_addr[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[4]~4 (
	.dataa(\MonAReg[6]~q ),
	.datab(address_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.cout());
defparam \ociram_addr[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_addr[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[5]~5 (
	.dataa(\MonAReg[7]~q ),
	.datab(address_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.cout());
defparam \ociram_addr[5]~5 .lut_mask = 16'hAACC;
defparam \ociram_addr[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[6]~6 (
	.dataa(\MonAReg[8]~q ),
	.datab(address_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.cout());
defparam \ociram_addr[6]~6 .lut_mask = 16'hAACC;
defparam \ociram_addr[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[7]~7 (
	.dataa(\MonAReg[9]~q ),
	.datab(address_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.cout());
defparam \ociram_addr[7]~7 .lut_mask = 16'hAACC;
defparam \ociram_addr[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.cout());
defparam \ociram_byteenable[0]~0 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(MonDReg_1),
	.datab(writedata_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.cout());
defparam \ociram_wr_data[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_wr~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_ram_wr~q ),
	.datac(jdo_35),
	.datad(\MonARegAddrInc[8]~16_combout ),
	.cin(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.cout());
defparam \jtag_ram_wr~0 .lut_mask = 16'hACFF;
defparam \jtag_ram_wr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(MonDReg_2),
	.datab(writedata_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.cout());
defparam \ociram_wr_data[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[3]~3 (
	.dataa(MonDReg_3),
	.datab(writedata_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[3]~3_combout ),
	.cout());
defparam \ociram_wr_data[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[4]~4 (
	.dataa(MonDReg_4),
	.datab(writedata_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[4]~4_combout ),
	.cout());
defparam \ociram_wr_data[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[21]~5 (
	.dataa(MonDReg_21),
	.datab(writedata_21),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[21]~5_combout ),
	.cout());
defparam \ociram_wr_data[21]~5 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[21]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.cout());
defparam \ociram_byteenable[2]~1 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[22]~6 (
	.dataa(MonDReg_22),
	.datab(writedata_22),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[22]~6_combout ),
	.cout());
defparam \ociram_wr_data[22]~6 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[22]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[23]~7 (
	.dataa(MonDReg_23),
	.datab(writedata_23),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[23]~7_combout ),
	.cout());
defparam \ociram_wr_data[23]~7 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[23]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[24]~8 (
	.dataa(MonDReg_24),
	.datab(writedata_24),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[24]~8_combout ),
	.cout());
defparam \ociram_wr_data[24]~8 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[24]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.cout());
defparam \ociram_byteenable[3]~2 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[25]~9 (
	.dataa(MonDReg_25),
	.datab(writedata_25),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[25]~9_combout ),
	.cout());
defparam \ociram_wr_data[25]~9 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[25]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[26]~10 (
	.dataa(MonDReg_26),
	.datab(writedata_26),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[26]~10_combout ),
	.cout());
defparam \ociram_wr_data[26]~10 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[26]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[11]~11 (
	.dataa(MonDReg_11),
	.datab(writedata_11),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[11]~11_combout ),
	.cout());
defparam \ociram_wr_data[11]~11 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[11]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.cout());
defparam \ociram_byteenable[1]~3 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[13]~12 (
	.dataa(MonDReg_13),
	.datab(writedata_13),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[13]~12_combout ),
	.cout());
defparam \ociram_wr_data[13]~12 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[13]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[16]~13 (
	.dataa(MonDReg_16),
	.datab(writedata_16),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[16]~13_combout ),
	.cout());
defparam \ociram_wr_data[16]~13 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[16]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[12]~14 (
	.dataa(MonDReg_12),
	.datab(writedata_12),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[12]~14_combout ),
	.cout());
defparam \ociram_wr_data[12]~14 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[12]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[5]~15 (
	.dataa(MonDReg_5),
	.datab(writedata_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[5]~15_combout ),
	.cout());
defparam \ociram_wr_data[5]~15 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[5]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[14]~16 (
	.dataa(MonDReg_14),
	.datab(writedata_14),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[14]~16_combout ),
	.cout());
defparam \ociram_wr_data[14]~16 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[14]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[15]~17 (
	.dataa(MonDReg_15),
	.datab(writedata_15),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[15]~17_combout ),
	.cout());
defparam \ociram_wr_data[15]~17 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[15]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[10]~18 (
	.dataa(MonDReg_10),
	.datab(writedata_10),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[10]~18_combout ),
	.cout());
defparam \ociram_wr_data[10]~18 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[10]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[9]~19 (
	.dataa(MonDReg_9),
	.datab(writedata_9),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[9]~19_combout ),
	.cout());
defparam \ociram_wr_data[9]~19 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[9]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[8]~20 (
	.dataa(MonDReg_8),
	.datab(writedata_8),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[8]~20_combout ),
	.cout());
defparam \ociram_wr_data[8]~20 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[8]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[7]~21 (
	.dataa(MonDReg_7),
	.datab(writedata_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[7]~21_combout ),
	.cout());
defparam \ociram_wr_data[7]~21 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[7]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[6]~22 (
	.dataa(MonDReg_6),
	.datab(writedata_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[6]~22_combout ),
	.cout());
defparam \ociram_wr_data[6]~22 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[6]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[20]~23 (
	.dataa(MonDReg_20),
	.datab(writedata_20),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[20]~23_combout ),
	.cout());
defparam \ociram_wr_data[20]~23 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[20]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[18]~24 (
	.dataa(MonDReg_18),
	.datab(writedata_18),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[18]~24_combout ),
	.cout());
defparam \ociram_wr_data[18]~24 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[18]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[19]~25 (
	.dataa(MonDReg_19),
	.datab(writedata_19),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[19]~25_combout ),
	.cout());
defparam \ociram_wr_data[19]~25 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[19]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[17]~26 (
	.dataa(MonDReg_17),
	.datab(writedata_17),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[17]~26_combout ),
	.cout());
defparam \ociram_wr_data[17]~26 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[17]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[27]~27 (
	.dataa(MonDReg_27),
	.datab(writedata_27),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[27]~27_combout ),
	.cout());
defparam \ociram_wr_data[27]~27 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[27]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[28]~28 (
	.dataa(MonDReg_28),
	.datab(writedata_28),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[28]~28_combout ),
	.cout());
defparam \ociram_wr_data[28]~28 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[28]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[31]~29 (
	.dataa(MonDReg_31),
	.datab(writedata_31),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[31]~29_combout ),
	.cout());
defparam \ociram_wr_data[31]~29 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[31]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[30]~30 (
	.dataa(MonDReg_30),
	.datab(writedata_30),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[30]~30_combout ),
	.cout());
defparam \ociram_wr_data[30]~30 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[30]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[29]~31 (
	.dataa(MonDReg_29),
	.datab(writedata_29),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[29]~31_combout ),
	.cout());
defparam \ociram_wr_data[29]~31 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[29]~31 .sum_lutc_input = "datac";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg[0]~0_combout ),
	.asdata(jdo_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg[2]~1_combout ),
	.asdata(jdo_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg[3]~2_combout ),
	.asdata(jdo_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg[4]~3_combout ),
	.asdata(jdo_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(\MonDReg[27]~4_combout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[27]~21_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg[11]~6_combout ),
	.asdata(jdo_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg[12]~7_combout ),
	.asdata(jdo_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg[5]~5_combout ),
	.asdata(jdo_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(\MonDReg[10]~11_combout ),
	.asdata(jdo_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~10_combout ),
	.asdata(jdo_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[27]~21_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg[18]~8_combout ),
	.asdata(jdo_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg[29]~9_combout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

cycloneive_lcell_comb \ociram_wr_en~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(ociram_wr_en),
	.cout());
defparam \ociram_wr_en~0 .lut_mask = 16'hEEEE;
defparam \ociram_wr_en~0 .sum_lutc_input = "datac";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(\MonDReg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(\MonDReg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(\MonDReg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(\MonDReg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(\MonDReg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(\MonDReg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(\MonDReg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(\MonDReg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(\MonDReg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(\MonDReg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(\MonDReg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(\MonDReg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(\MonDReg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(\MonDReg~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\MonARegAddrInc[0]~0_combout ),
	.cout(\MonARegAddrInc[0]~1 ));
defparam \MonARegAddrInc[0]~0 .lut_mask = 16'h55AA;
defparam \MonARegAddrInc[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonAReg~0 (
	.dataa(\MonARegAddrInc[0]~0_combout ),
	.datab(jdo_26),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~0_combout ),
	.cout());
defparam \MonAReg~0 .lut_mask = 16'hAACC;
defparam \MonAReg~0 .sum_lutc_input = "datac";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\MonAReg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[1]~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[0]~1 ),
	.combout(\MonARegAddrInc[1]~2_combout ),
	.cout(\MonARegAddrInc[1]~3 ));
defparam \MonARegAddrInc[1]~2 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~2 (
	.dataa(\MonARegAddrInc[1]~2_combout ),
	.datab(jdo_27),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~2_combout ),
	.cout());
defparam \MonAReg~2 .lut_mask = 16'hAACC;
defparam \MonAReg~2 .sum_lutc_input = "datac";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\MonAReg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[2]~4 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[1]~3 ),
	.combout(\MonARegAddrInc[2]~4_combout ),
	.cout(\MonARegAddrInc[2]~5 ));
defparam \MonARegAddrInc[2]~4 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~1 (
	.dataa(\MonARegAddrInc[2]~4_combout ),
	.datab(jdo_28),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~1_combout ),
	.cout());
defparam \MonAReg~1 .lut_mask = 16'hAACC;
defparam \MonAReg~1 .sum_lutc_input = "datac";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\MonAReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonAReg~3 (
	.dataa(\MonARegAddrInc[8]~16_combout ),
	.datab(jdo_17),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~3_combout ),
	.cout());
defparam \MonAReg~3 .lut_mask = 16'hAACC;
defparam \MonAReg~3 .sum_lutc_input = "datac";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\MonAReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[3]~6 (
	.dataa(\MonAReg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[2]~5 ),
	.combout(\MonARegAddrInc[3]~6_combout ),
	.cout(\MonARegAddrInc[3]~7 ));
defparam \MonARegAddrInc[3]~6 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~8 (
	.dataa(\MonARegAddrInc[3]~6_combout ),
	.datab(jdo_29),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~8_combout ),
	.cout());
defparam \MonAReg~8 .lut_mask = 16'hAACC;
defparam \MonAReg~8 .sum_lutc_input = "datac";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\MonAReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[4]~8 (
	.dataa(\MonAReg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[3]~7 ),
	.combout(\MonARegAddrInc[4]~8_combout ),
	.cout(\MonARegAddrInc[4]~9 ));
defparam \MonARegAddrInc[4]~8 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[4]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~7 (
	.dataa(\MonARegAddrInc[4]~8_combout ),
	.datab(jdo_30),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~7_combout ),
	.cout());
defparam \MonAReg~7 .lut_mask = 16'hAACC;
defparam \MonAReg~7 .sum_lutc_input = "datac";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\MonAReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[5]~10 (
	.dataa(\MonAReg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[4]~9 ),
	.combout(\MonARegAddrInc[5]~10_combout ),
	.cout(\MonARegAddrInc[5]~11 ));
defparam \MonARegAddrInc[5]~10 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~6 (
	.dataa(\MonARegAddrInc[5]~10_combout ),
	.datab(jdo_31),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~6_combout ),
	.cout());
defparam \MonAReg~6 .lut_mask = 16'hAACC;
defparam \MonAReg~6 .sum_lutc_input = "datac";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\MonAReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[6]~12 (
	.dataa(\MonAReg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[5]~11 ),
	.combout(\MonARegAddrInc[6]~12_combout ),
	.cout(\MonARegAddrInc[6]~13 ));
defparam \MonARegAddrInc[6]~12 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~5 (
	.dataa(\MonARegAddrInc[6]~12_combout ),
	.datab(jdo_32),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~5_combout ),
	.cout());
defparam \MonAReg~5 .lut_mask = 16'hAACC;
defparam \MonAReg~5 .sum_lutc_input = "datac";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\MonAReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[7]~14 (
	.dataa(\MonAReg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[6]~13 ),
	.combout(\MonARegAddrInc[7]~14_combout ),
	.cout(\MonARegAddrInc[7]~15 ));
defparam \MonARegAddrInc[7]~14 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~4 (
	.dataa(\MonARegAddrInc[7]~14_combout ),
	.datab(jdo_33),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~4_combout ),
	.cout());
defparam \MonAReg~4 .lut_mask = 16'hAACC;
defparam \MonAReg~4 .sum_lutc_input = "datac";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\MonAReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[8]~16 (
	.dataa(\MonAReg[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\MonARegAddrInc[7]~15 ),
	.combout(\MonARegAddrInc[8]~16_combout ),
	.cout());
defparam \MonARegAddrInc[8]~16 .lut_mask = 16'h5A5A;
defparam \MonARegAddrInc[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \jtag_ram_rd~0 (
	.dataa(jdo_35),
	.datab(\jtag_ram_rd~q ),
	.datac(jdo_34),
	.datad(\MonARegAddrInc[8]~16_combout ),
	.cin(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.cout());
defparam \jtag_ram_rd~0 .lut_mask = 16'hF7B3;
defparam \jtag_ram_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_rd~1 (
	.dataa(take_action_ocimem_a),
	.datab(take_action_ocimem_a1),
	.datac(jdo_17),
	.datad(\jtag_ram_rd~0_combout ),
	.cin(gnd),
	.combout(\jtag_ram_rd~1_combout ),
	.cout());
defparam \jtag_ram_rd~1 .lut_mask = 16'hEFFF;
defparam \jtag_ram_rd~1 .sum_lutc_input = "datac";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~0 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_0),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[0]~0_combout ),
	.cout());
defparam \MonDReg[0]~0 .lut_mask = 16'hAACC;
defparam \MonDReg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_rd~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_rd~q ),
	.datac(gnd),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\jtag_rd~0_combout ),
	.cout());
defparam \jtag_rd~0 .lut_mask = 16'hEEFF;
defparam \jtag_rd~0 .sum_lutc_input = "datac";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(\jtag_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~12 (
	.dataa(gnd),
	.datab(take_action_ocimem_a),
	.datac(\jtag_rd_d1~q ),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\MonDReg[0]~12_combout ),
	.cout());
defparam \MonDReg[0]~12 .lut_mask = 16'hF3C0;
defparam \MonDReg[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[2]~1 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_2),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[2]~1_combout ),
	.cout());
defparam \MonDReg[2]~1 .lut_mask = 16'hAACC;
defparam \MonDReg[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[3]~2 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_3),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[3]~2_combout ),
	.cout());
defparam \MonDReg[3]~2 .lut_mask = 16'hAACC;
defparam \MonDReg[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[4]~3 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_4),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[4]~3_combout ),
	.cout());
defparam \MonDReg[4]~3 .lut_mask = 16'hAACC;
defparam \MonDReg[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cfgrom_readdata[27]~0 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\cfgrom_readdata[27]~0_combout ),
	.cout());
defparam \cfgrom_readdata[27]~0 .lut_mask = 16'hAFFA;
defparam \cfgrom_readdata[27]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[27]~4 (
	.dataa(\cfgrom_readdata[27]~0_combout ),
	.datab(q_a_27),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[27]~4_combout ),
	.cout());
defparam \MonDReg[27]~4 .lut_mask = 16'hCC55;
defparam \MonDReg[27]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[27]~21 (
	.dataa(take_action_ocimem_b),
	.datab(\jtag_rd_d1~q ),
	.datac(gnd),
	.datad(take_action_ocimem_a),
	.cin(gnd),
	.combout(\MonDReg[27]~21_combout ),
	.cout());
defparam \MonDReg[27]~21 .lut_mask = 16'hEEFF;
defparam \MonDReg[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[11]~6 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_11),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[11]~6_combout ),
	.cout());
defparam \MonDReg[11]~6 .lut_mask = 16'hAACC;
defparam \MonDReg[11]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[12]~7 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_12),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[12]~7_combout ),
	.cout());
defparam \MonDReg[12]~7 .lut_mask = 16'hAACC;
defparam \MonDReg[12]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(gnd),
	.datab(\MonAReg[2]~q ),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h3FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[5]~5 (
	.dataa(\Equal0~1_combout ),
	.datab(q_a_5),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[5]~5_combout ),
	.cout());
defparam \MonDReg[5]~5 .lut_mask = 16'hAACC;
defparam \MonDReg[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[10]~11 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_10),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[10]~11_combout ),
	.cout());
defparam \MonDReg[10]~11 .lut_mask = 16'hAACC;
defparam \MonDReg[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cfgrom_readdata[8]~1 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\cfgrom_readdata[8]~1_combout ),
	.cout());
defparam \cfgrom_readdata[8]~1 .lut_mask = 16'hAAFF;
defparam \cfgrom_readdata[8]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[8]~10 (
	.dataa(\cfgrom_readdata[8]~1_combout ),
	.datab(q_a_8),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[8]~10_combout ),
	.cout());
defparam \MonDReg[8]~10 .lut_mask = 16'hAACC;
defparam \MonDReg[8]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hAFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[18]~8 (
	.dataa(\Equal0~2_combout ),
	.datab(q_a_18),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[18]~8_combout ),
	.cout());
defparam \MonDReg[18]~8 .lut_mask = 16'hAACC;
defparam \MonDReg[18]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hAFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[29]~9 (
	.dataa(\Equal0~3_combout ),
	.datab(q_a_29),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[29]~9_combout ),
	.cout());
defparam \MonDReg[29]~9 .lut_mask = 16'hAACC;
defparam \MonDReg[29]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~0 (
	.dataa(jdo_34),
	.datab(gnd),
	.datac(gnd),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.cout());
defparam \jtag_ram_access~0 .lut_mask = 16'hAAFF;
defparam \jtag_ram_access~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~1 (
	.dataa(jdo_17),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(\jtag_ram_access~0_combout ),
	.datad(take_action_ocimem_a),
	.cin(gnd),
	.combout(\jtag_ram_access~1_combout ),
	.cout());
defparam \jtag_ram_access~1 .lut_mask = 16'hF737;
defparam \jtag_ram_access~1 .sum_lutc_input = "datac";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cycloneive_lcell_comb \waitrequest~0 (
	.dataa(write),
	.datab(\jtag_ram_access~q ),
	.datac(address_8),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\waitrequest~0_combout ),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hEFFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(read),
	.datab(address_8),
	.datac(\jtag_ram_access~q ),
	.datad(write),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 16'hEFFF;
defparam \avalon_ociram_readdata_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~1 (
	.dataa(waitrequest1),
	.datab(\avalon_ociram_readdata_ready~0_combout ),
	.datac(write),
	.datad(\avalon_ociram_readdata_ready~q ),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~1_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~1 .lut_mask = 16'hFFFE;
defparam \avalon_ociram_readdata_ready~1 .sum_lutc_input = "datac";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cycloneive_lcell_comb \waitrequest~1 (
	.dataa(\waitrequest~0_combout ),
	.datab(read),
	.datac(\avalon_ociram_readdata_ready~q ),
	.datad(write),
	.cin(gnd),
	.combout(\waitrequest~1_combout ),
	.cout());
defparam \waitrequest~1 .lut_mask = 16'hBFFF;
defparam \waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~13 (
	.dataa(jdo_4),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_1),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~13_combout ),
	.cout());
defparam \MonDReg~13 .lut_mask = 16'hFAFC;
defparam \MonDReg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~14 (
	.dataa(jdo_24),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_21),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~14_combout ),
	.cout());
defparam \MonDReg~14 .lut_mask = 16'hFAFC;
defparam \MonDReg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~15 (
	.dataa(jdo_25),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_22),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~15_combout ),
	.cout());
defparam \MonDReg~15 .lut_mask = 16'hFAFC;
defparam \MonDReg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~16 (
	.dataa(jdo_19),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_16),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~16_combout ),
	.cout());
defparam \MonDReg~16 .lut_mask = 16'hFAFC;
defparam \MonDReg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~17 (
	.dataa(jdo_23),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_20),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~17_combout ),
	.cout());
defparam \MonDReg~17 .lut_mask = 16'hFAFC;
defparam \MonDReg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~18 (
	.dataa(jdo_22),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_19),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~18_combout ),
	.cout());
defparam \MonDReg~18 .lut_mask = 16'hFAFC;
defparam \MonDReg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~19 (
	.dataa(jdo_26),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_23),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~19_combout ),
	.cout());
defparam \MonDReg~19 .lut_mask = 16'hFAFC;
defparam \MonDReg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~20 (
	.dataa(jdo_28),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_25),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~20_combout ),
	.cout());
defparam \MonDReg~20 .lut_mask = 16'hFAFC;
defparam \MonDReg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~22 (
	.dataa(jdo_29),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_26),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~22_combout ),
	.cout());
defparam \MonDReg~22 .lut_mask = 16'hFAFC;
defparam \MonDReg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~23 (
	.dataa(jdo_27),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_24),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~23_combout ),
	.cout());
defparam \MonDReg~23 .lut_mask = 16'hFAFC;
defparam \MonDReg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~24 (
	.dataa(jdo_16),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_13),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~24_combout ),
	.cout());
defparam \MonDReg~24 .lut_mask = 16'hFAFC;
defparam \MonDReg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~25 (
	.dataa(jdo_17),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_14),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~25_combout ),
	.cout());
defparam \MonDReg~25 .lut_mask = 16'hFAFC;
defparam \MonDReg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~26 (
	.dataa(jdo_18),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_15),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~26_combout ),
	.cout());
defparam \MonDReg~26 .lut_mask = 16'hFAFC;
defparam \MonDReg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~27 (
	.dataa(jdo_12),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_9),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~27_combout ),
	.cout());
defparam \MonDReg~27 .lut_mask = 16'hFAFC;
defparam \MonDReg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~28 (
	.dataa(jdo_10),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_7),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~28_combout ),
	.cout());
defparam \MonDReg~28 .lut_mask = 16'hFAFC;
defparam \MonDReg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~29 (
	.dataa(jdo_9),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_6),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~29_combout ),
	.cout());
defparam \MonDReg~29 .lut_mask = 16'hFAFC;
defparam \MonDReg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~30 (
	.dataa(jdo_20),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_17),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~30_combout ),
	.cout());
defparam \MonDReg~30 .lut_mask = 16'hFAFC;
defparam \MonDReg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~31 (
	.dataa(jdo_31),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_28),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~31_combout ),
	.cout());
defparam \MonDReg~31 .lut_mask = 16'hFAFC;
defparam \MonDReg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~32 (
	.dataa(jdo_34),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_31),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~32_combout ),
	.cout());
defparam \MonDReg~32 .lut_mask = 16'hFAFC;
defparam \MonDReg~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~33 (
	.dataa(jdo_33),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_30),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~33_combout ),
	.cout());
defparam \MonDReg~33 .lut_mask = 16'hFAFC;
defparam \MonDReg~33 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_cpu_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_21,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_18,
	q_a_19,
	q_a_17,
	q_a_27,
	q_a_28,
	q_a_31,
	q_a_30,
	q_a_29,
	ociram_wr_en,
	r_early_rst,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_3,
	ociram_wr_data_4,
	ociram_wr_data_21,
	ociram_byteenable_2,
	ociram_wr_data_22,
	ociram_wr_data_23,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_25,
	ociram_wr_data_26,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_13,
	ociram_wr_data_16,
	ociram_wr_data_12,
	ociram_wr_data_5,
	ociram_wr_data_14,
	ociram_wr_data_15,
	ociram_wr_data_10,
	ociram_wr_data_9,
	ociram_wr_data_8,
	ociram_wr_data_7,
	ociram_wr_data_6,
	ociram_wr_data_20,
	ociram_wr_data_18,
	ociram_wr_data_19,
	ociram_wr_data_17,
	ociram_wr_data_27,
	ociram_wr_data_28,
	ociram_wr_data_31,
	ociram_wr_data_30,
	ociram_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_21;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_18;
output 	q_a_19;
output 	q_a_17;
output 	q_a_27;
output 	q_a_28;
output 	q_a_31;
output 	q_a_30;
output 	q_a_29;
input 	ociram_wr_en;
input 	r_early_rst;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_3;
input 	ociram_wr_data_4;
input 	ociram_wr_data_21;
input 	ociram_byteenable_2;
input 	ociram_wr_data_22;
input 	ociram_wr_data_23;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_25;
input 	ociram_wr_data_26;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_13;
input 	ociram_wr_data_16;
input 	ociram_wr_data_12;
input 	ociram_wr_data_5;
input 	ociram_wr_data_14;
input 	ociram_wr_data_15;
input 	ociram_wr_data_10;
input 	ociram_wr_data_9;
input 	ociram_wr_data_8;
input 	ociram_wr_data_7;
input 	ociram_wr_data_6;
input 	ociram_wr_data_20;
input 	ociram_wr_data_18;
input 	ociram_wr_data_19;
input 	ociram_wr_data_17;
input 	ociram_wr_data_27;
input 	ociram_wr_data_28;
input 	ociram_wr_data_31;
input 	ociram_wr_data_30;
input 	ociram_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(r_early_rst),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module usb_system_altsyncram_1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_4a31 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module usb_system_altsyncram_4a31 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_nios2_oci:the_usb_system_cpu_cpu_nios2_oci|usb_system_cpu_cpu_nios2_ocimem:the_usb_system_cpu_cpu_nios2_ocimem|usb_system_cpu_cpu_ociram_sp_ram_module:usb_system_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module usb_system_usb_system_cpu_cpu_register_bank_a_module (
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_24,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_31,
	q_b_29,
	q_b_30,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	D_iw_27,
	D_iw_28,
	D_iw_31,
	D_iw_30,
	D_iw_29,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_8,
	W_rf_wr_data_9,
	W_rf_wr_data_10,
	W_rf_wr_data_11,
	W_rf_wr_data_12,
	W_rf_wr_data_13,
	W_rf_wr_data_14,
	W_rf_wr_data_15,
	W_rf_wr_data_16,
	W_rf_wr_data_17,
	W_rf_wr_data_18,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_24,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_31,
	W_rf_wr_data_29,
	W_rf_wr_data_30,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_24;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_31;
output 	q_b_29;
output 	q_b_30;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	D_iw_27;
input 	D_iw_28;
input 	D_iw_31;
input 	D_iw_30;
input 	D_iw_29;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_30;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.address_b({D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.clock0(clk_clk));

endmodule

module usb_system_altsyncram_2 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_6mc1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module usb_system_altsyncram_6mc1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_a_module:usb_system_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

endmodule

module usb_system_usb_system_cpu_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_24,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_31,
	q_b_29,
	q_b_30,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	D_iw_22,
	D_iw_23,
	D_iw_24,
	D_iw_25,
	D_iw_26,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_8,
	W_rf_wr_data_9,
	W_rf_wr_data_10,
	W_rf_wr_data_11,
	W_rf_wr_data_12,
	W_rf_wr_data_13,
	W_rf_wr_data_14,
	W_rf_wr_data_15,
	W_rf_wr_data_16,
	W_rf_wr_data_17,
	W_rf_wr_data_18,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_24,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_31,
	W_rf_wr_data_29,
	W_rf_wr_data_30,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_24;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_31;
output 	q_b_29;
output 	q_b_30;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	D_iw_22;
input 	D_iw_23;
input 	D_iw_24;
input 	D_iw_25;
input 	D_iw_26;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_30;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_3 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.address_b({D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.clock0(clk_clk));

endmodule

module usb_system_altsyncram_3 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_6mc1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module usb_system_altsyncram_6mc1_1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "usb_system_cpu:cpu|usb_system_cpu_cpu:cpu|usb_system_cpu_cpu_register_bank_b_module:usb_system_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

endmodule

module usb_system_usb_system_jtag_uart (
	W_alu_result_2,
	tdo,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_10,
	sink_in_reset,
	d_read,
	read_accepted,
	uav_write,
	mem_used_1,
	av_waitrequest1,
	Equal9,
	s0_cmd_valid,
	sink_ready,
	av_readdata_9,
	av_readdata_8,
	b_full,
	read_01,
	av_readdata_0,
	av_readdata_1,
	av_readdata_2,
	av_readdata_3,
	av_readdata_4,
	av_readdata_5,
	av_readdata_6,
	av_readdata_7,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_01,
	counter_reg_bit_11,
	counter_reg_bit_41,
	counter_reg_bit_51,
	ac1,
	woverflow1,
	rvalid1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
output 	tdo;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_10;
input 	sink_in_reset;
input 	d_read;
input 	read_accepted;
input 	uav_write;
input 	mem_used_1;
output 	av_waitrequest1;
input 	Equal9;
input 	s0_cmd_valid;
input 	sink_ready;
output 	av_readdata_9;
output 	av_readdata_8;
output 	b_full;
output 	read_01;
output 	av_readdata_0;
output 	av_readdata_1;
output 	av_readdata_2;
output 	av_readdata_3;
output 	av_readdata_4;
output 	av_readdata_5;
output 	av_readdata_6;
output 	av_readdata_7;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	counter_reg_bit_31;
output 	counter_reg_bit_21;
output 	counter_reg_bit_01;
output 	counter_reg_bit_11;
output 	counter_reg_bit_41;
output 	counter_reg_bit_51;
output 	ac1;
output 	woverflow1;
output 	rvalid1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ;
wire \the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ;
wire \t_dav~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|r_ena1~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|t_pause~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|t_ena~q ;
wire \the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_wr~q ;
wire \wr_rfifo~combout ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[0]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[1]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[2]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[3]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[4]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[5]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[6]~q ;
wire \usb_system_jtag_uart_alt_jtag_atlantic|wdata[7]~q ;
wire \fifo_wr~0_combout ;
wire \always2~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \fifo_rd~0_combout ;
wire \ien_AF~0_combout ;
wire \ien_AE~q ;
wire \ien_AF~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~0_combout ;
wire \Add0~2_combout ;
wire \LessThan1~0_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \LessThan1~1_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \LessThan1~2_combout ;
wire \fifo_AF~q ;
wire \fifo_rd~1_combout ;
wire \fifo_rd~2_combout ;
wire \ac~0_combout ;
wire \ac~1_combout ;
wire \woverflow~0_combout ;
wire \woverflow~1_combout ;
wire \rvalid~0_combout ;
wire \rvalid~1_combout ;


usb_system_usb_system_jtag_uart_scfifo_r the_usb_system_jtag_uart_scfifo_r(
	.q_b_0(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ),
	.q_b_1(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ),
	.q_b_2(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ),
	.q_b_3(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ),
	.q_b_4(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ),
	.q_b_5(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ),
	.q_b_6(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ),
	.q_b_7(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_31),
	.counter_reg_bit_2(counter_reg_bit_21),
	.counter_reg_bit_0(counter_reg_bit_01),
	.counter_reg_bit_1(counter_reg_bit_11),
	.counter_reg_bit_4(counter_reg_bit_41),
	.counter_reg_bit_5(counter_reg_bit_51),
	.t_ena(\usb_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.rvalid(\rvalid~0_combout ),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.clk_clk(clk_clk));

usb_system_usb_system_jtag_uart_scfifo_w the_usb_system_jtag_uart_scfifo_w(
	.q_b_7(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ),
	.q_b_0(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ),
	.q_b_1(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ),
	.q_b_2(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ),
	.q_b_3(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ),
	.q_b_4(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ),
	.q_b_5(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ),
	.q_b_6(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.fifo_wr(\fifo_wr~q ),
	.clk_clk(clk_clk));

usb_system_alt_jtag_atlantic usb_system_jtag_uart_alt_jtag_atlantic(
	.r_dat({\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ,\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ,
\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ,\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ,
\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ,\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ,
\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ,\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] }),
	.tdo1(tdo),
	.rst_n(r_sync_rst),
	.sink_in_reset(sink_in_reset),
	.t_dav(\t_dav~q ),
	.rvalid01(\usb_system_jtag_uart_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\usb_system_jtag_uart_alt_jtag_atlantic|r_ena1~q ),
	.t_pause1(\usb_system_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.t_ena1(\usb_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.wdata_0(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\usb_system_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

cycloneive_lcell_comb \r_val~0 (
	.dataa(\the_usb_system_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datab(\r_val~q ),
	.datac(\usb_system_jtag_uart_alt_jtag_atlantic|r_ena1~q ),
	.datad(\usb_system_jtag_uart_alt_jtag_atlantic|rvalid0~q ),
	.cin(gnd),
	.combout(\r_val~0_combout ),
	.cout());
defparam \r_val~0 .lut_mask = 16'hBFFF;
defparam \r_val~0 .sum_lutc_input = "datac";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cycloneive_lcell_comb wr_rfifo(
	.dataa(\usb_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(b_full),
	.cin(gnd),
	.combout(\wr_rfifo~combout ),
	.cout());
defparam wr_rfifo.lut_mask = 16'hAAFF;
defparam wr_rfifo.sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_wr~0 (
	.dataa(W_alu_result_2),
	.datab(b_full1),
	.datac(uav_write),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\fifo_wr~0_combout ),
	.cout());
defparam \fifo_wr~0 .lut_mask = 16'hFFF7;
defparam \fifo_wr~0 .sum_lutc_input = "datac";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

cycloneive_lcell_comb \av_readdata[9] (
	.dataa(\fifo_AE~q ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_9),
	.cout());
defparam \av_readdata[9] .lut_mask = 16'hEEEE;
defparam \av_readdata[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[8]~0 (
	.dataa(\ien_AF~q ),
	.datab(\pause_irq~q ),
	.datac(\fifo_AF~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_8),
	.cout());
defparam \av_readdata[8]~0 .lut_mask = 16'hFEFE;
defparam \av_readdata[8]~0 .sum_lutc_input = "datac";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

cycloneive_lcell_comb \av_readdata[0]~1 (
	.dataa(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ),
	.datab(\ien_AF~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_0),
	.cout());
defparam \av_readdata[0]~1 .lut_mask = 16'hAACC;
defparam \av_readdata[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[1]~2 (
	.dataa(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_1),
	.cout());
defparam \av_readdata[1]~2 .lut_mask = 16'hAACC;
defparam \av_readdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[2]~3 (
	.dataa(read_01),
	.datab(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_2),
	.cout());
defparam \av_readdata[2]~3 .lut_mask = 16'hEEEE;
defparam \av_readdata[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[3]~4 (
	.dataa(read_01),
	.datab(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_3),
	.cout());
defparam \av_readdata[3]~4 .lut_mask = 16'hEEEE;
defparam \av_readdata[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[4]~5 (
	.dataa(read_01),
	.datab(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_4),
	.cout());
defparam \av_readdata[4]~5 .lut_mask = 16'hEEEE;
defparam \av_readdata[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[5]~6 (
	.dataa(read_01),
	.datab(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_5),
	.cout());
defparam \av_readdata[5]~6 .lut_mask = 16'hEEEE;
defparam \av_readdata[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[6]~7 (
	.dataa(read_01),
	.datab(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_6),
	.cout());
defparam \av_readdata[6]~7 .lut_mask = 16'hEEEE;
defparam \av_readdata[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[7]~8 (
	.dataa(read_01),
	.datab(\the_usb_system_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_7),
	.cout());
defparam \av_readdata[7]~8 .lut_mask = 16'hEEEE;
defparam \av_readdata[7]~8 .sum_lutc_input = "datac";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cycloneive_lcell_comb \always2~0 (
	.dataa(Equal9),
	.datab(s0_cmd_valid),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hEFFF;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hFFFE;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\LessThan0~0_combout ),
	.datab(b_full1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cycloneive_lcell_comb \fifo_rd~0 (
	.dataa(Equal9),
	.datab(gnd),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\fifo_rd~0_combout ),
	.cout());
defparam \fifo_rd~0 .lut_mask = 16'hAFFF;
defparam \fifo_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ien_AF~0 (
	.dataa(W_alu_result_2),
	.datab(uav_write),
	.datac(s0_cmd_valid),
	.datad(\fifo_rd~0_combout ),
	.cin(gnd),
	.combout(\ien_AF~0_combout ),
	.cout());
defparam \ien_AF~0 .lut_mask = 16'hFFFE;
defparam \ien_AF~0 .sum_lutc_input = "datac";

dffeas ien_AE(
	.clk(clk_clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~0_combout ),
	.q(\ien_AE~q ),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

dffeas ien_AF(
	.clk(clk_clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~0_combout ),
	.q(\ien_AF~q ),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cycloneive_lcell_comb \pause_irq~0 (
	.dataa(b_non_empty),
	.datab(\usb_system_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.datac(\pause_irq~q ),
	.datad(read_01),
	.cin(gnd),
	.combout(\pause_irq~0_combout ),
	.cout());
defparam \pause_irq~0 .lut_mask = 16'hFEFF;
defparam \pause_irq~0 .sum_lutc_input = "datac";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(counter_reg_bit_01),
	.datab(counter_reg_bit_11),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h6677;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~2 (
	.dataa(counter_reg_bit_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5AAF;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(counter_reg_bit_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5A5F;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~0 (
	.dataa(\Add0~4_combout ),
	.datab(counter_reg_bit_01),
	.datac(\Add0~0_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hFFFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~6 (
	.dataa(counter_reg_bit_41),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5AAF;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~8 (
	.dataa(counter_reg_bit_51),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~1 (
	.dataa(\Add0~6_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
defparam \LessThan1~1 .lut_mask = 16'hEEEE;
defparam \LessThan1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~10 (
	.dataa(b_full),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5AAF;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'hF0F0;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~2 (
	.dataa(\LessThan1~0_combout ),
	.datab(\LessThan1~1_combout ),
	.datac(\Add0~10_combout ),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\LessThan1~2_combout ),
	.cout());
defparam \LessThan1~2 .lut_mask = 16'h7FFF;
defparam \LessThan1~2 .sum_lutc_input = "datac";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cycloneive_lcell_comb \fifo_rd~1 (
	.dataa(d_read),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(read_accepted),
	.cin(gnd),
	.combout(\fifo_rd~1_combout ),
	.cout());
defparam \fifo_rd~1 .lut_mask = 16'hAFFF;
defparam \fifo_rd~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_rd~2 (
	.dataa(Equal9),
	.datab(\fifo_rd~1_combout ),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\fifo_rd~2_combout ),
	.cout());
defparam \fifo_rd~2 .lut_mask = 16'hEFFF;
defparam \fifo_rd~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~0 (
	.dataa(\usb_system_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.datab(\usb_system_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac~0_combout ),
	.cout());
defparam \ac~0 .lut_mask = 16'hEEEE;
defparam \ac~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~1 (
	.dataa(\ac~0_combout ),
	.datab(ac1),
	.datac(d_writedata_10),
	.datad(\ien_AF~0_combout ),
	.cin(gnd),
	.combout(\ac~1_combout ),
	.cout());
defparam \ac~1 .lut_mask = 16'hEFFF;
defparam \ac~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~0 (
	.dataa(uav_write),
	.datab(s0_cmd_valid),
	.datac(\fifo_rd~0_combout ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\woverflow~0_combout ),
	.cout());
defparam \woverflow~0 .lut_mask = 16'hFEFF;
defparam \woverflow~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~1 (
	.dataa(b_full1),
	.datab(woverflow1),
	.datac(gnd),
	.datad(\woverflow~0_combout ),
	.cin(gnd),
	.combout(\woverflow~1_combout ),
	.cout());
defparam \woverflow~1 .lut_mask = 16'hAACC;
defparam \woverflow~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rvalid~0 (
	.dataa(sink_ready),
	.datab(b_non_empty),
	.datac(\fifo_rd~1_combout ),
	.datad(av_waitrequest1),
	.cin(gnd),
	.combout(\rvalid~0_combout ),
	.cout());
defparam \rvalid~0 .lut_mask = 16'hFEFF;
defparam \rvalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rvalid~1 (
	.dataa(\rvalid~0_combout ),
	.datab(rvalid1),
	.datac(\fifo_rd~0_combout ),
	.datad(\fifo_rd~1_combout ),
	.cin(gnd),
	.combout(\rvalid~1_combout ),
	.cout());
defparam \rvalid~1 .lut_mask = 16'hEFFF;
defparam \rvalid~1 .sum_lutc_input = "datac";

endmodule

module usb_system_alt_jtag_atlantic (
	r_dat,
	tdo1,
	rst_n,
	sink_in_reset,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_pause1,
	t_ena1,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	tdo1;
input 	rst_n;
input 	sink_in_reset;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_pause1;
output 	t_ena1;
output 	wdata_0;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	wdata_6;
output 	wdata_7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \count~2_combout ;
wire \td_shift[0]~4_combout ;
wire \count[1]~q ;
wire \count~10_combout ;
wire \count[2]~q ;
wire \count~9_combout ;
wire \count[3]~q ;
wire \count~8_combout ;
wire \count[4]~q ;
wire \count~7_combout ;
wire \count[5]~q ;
wire \count~6_combout ;
wire \count[6]~q ;
wire \count~5_combout ;
wire \count[7]~q ;
wire \count~3_combout ;
wire \count[8]~q ;
wire \always0~0_combout ;
wire \state~0_combout ;
wire \state~1_combout ;
wire \state~2_combout ;
wire \state~q ;
wire \count[9]~0_combout ;
wire \count[9]~1_combout ;
wire \count[9]~q ;
wire \count~4_combout ;
wire \count[0]~q ;
wire \wdata[1]~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~1_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift~11_combout ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~8_combout ;
wire \td_shift[9]~q ;
wire \td_shift~6_combout ;
wire \rdata[6]~q ;
wire \td_shift~22_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~20_combout ;
wire \td_shift~21_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~18_combout ;
wire \td_shift~19_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~16_combout ;
wire \td_shift~17_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~14_combout ;
wire \td_shift~15_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~12_combout ;
wire \td_shift~13_combout ;
wire \td_shift[3]~q ;
wire \rdata[0]~q ;
wire \td_shift~9_combout ;
wire \td_shift~10_combout ;
wire \td_shift[2]~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~2_combout ;
wire \write_stalled~q ;
wire \td_shift~5_combout ;
wire \td_shift~7_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~0_combout ;
wire \td_shift~1_combout ;
wire \td_shift~2_combout ;
wire \td_shift~3_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \read_req~q ;
wire \rvalid0~1_combout ;
wire \rst2~q ;
wire \rvalid0~2_combout ;
wire \write~0_combout ;
wire \wdata[1]~1_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~0_combout ;
wire \write_valid~q ;
wire \t_pause~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \t_pause~1_combout ;
wire \t_ena~2_combout ;
wire \t_ena~3_combout ;


dffeas tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tdo1),
	.prn(vcc));
defparam tdo.is_wysiwyg = "true";
defparam tdo.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~2_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas t_pause(
	.clk(clk),
	.d(\t_pause~1_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause1),
	.prn(vcc));
defparam t_pause.is_wysiwyg = "true";
defparam t_pause.power_up = "low";

dffeas t_ena(
	.clk(clk),
	.d(\t_ena~3_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena1),
	.prn(vcc));
defparam t_ena.is_wysiwyg = "true";
defparam t_ena.power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

cycloneive_lcell_comb \tck_t_dav~0 (
	.dataa(t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tck_t_dav~0_combout ),
	.cout());
defparam \tck_t_dav~0 .lut_mask = 16'h5555;
defparam \tck_t_dav~0 .sum_lutc_input = "datac";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cycloneive_lcell_comb \count~2 (
	.dataa(state_4),
	.datab(\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~2_combout ),
	.cout());
defparam \count~2 .lut_mask = 16'hEEEE;
defparam \count~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift[0]~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(state_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\td_shift[0]~4_combout ),
	.cout());
defparam \td_shift[0]~4 .lut_mask = 16'hFEFF;
defparam \td_shift[0]~4 .sum_lutc_input = "datac";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \count~10 (
	.dataa(\count[1]~q ),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~10_combout ),
	.cout());
defparam \count~10 .lut_mask = 16'hEEEE;
defparam \count~10 .sum_lutc_input = "datac";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count~9 (
	.dataa(state_4),
	.datab(\count[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~9_combout ),
	.cout());
defparam \count~9 .lut_mask = 16'hEEEE;
defparam \count~9 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count~8 (
	.dataa(state_4),
	.datab(\count[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~8_combout ),
	.cout());
defparam \count~8 .lut_mask = 16'hEEEE;
defparam \count~8 .sum_lutc_input = "datac";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count~7 (
	.dataa(state_4),
	.datab(\count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~7_combout ),
	.cout());
defparam \count~7 .lut_mask = 16'hEEEE;
defparam \count~7 .sum_lutc_input = "datac";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count~6 (
	.dataa(state_4),
	.datab(\count[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~6_combout ),
	.cout());
defparam \count~6 .lut_mask = 16'hEEEE;
defparam \count~6 .sum_lutc_input = "datac";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count~5 (
	.dataa(state_4),
	.datab(\count[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEEEE;
defparam \count~5 .sum_lutc_input = "datac";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \count~3 (
	.dataa(state_4),
	.datab(\count[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hEEEE;
defparam \count~3 .sum_lutc_input = "datac";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(gnd),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~0 (
	.dataa(state_4),
	.datab(\always0~0_combout ),
	.datac(altera_internal_jtag1),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hFEFF;
defparam \state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~1 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'h7777;
defparam \state~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~2 (
	.dataa(\state~q ),
	.datab(virtual_ir_scan_reg),
	.datac(\state~0_combout ),
	.datad(\state~1_combout ),
	.cin(gnd),
	.combout(\state~2_combout ),
	.cout());
defparam \state~2 .lut_mask = 16'hFFD8;
defparam \state~2 .sum_lutc_input = "datac";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cycloneive_lcell_comb \count[9]~0 (
	.dataa(altera_internal_jtag1),
	.datab(irf_reg_0_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[9]~0_combout ),
	.cout());
defparam \count[9]~0 .lut_mask = 16'hBBBB;
defparam \count[9]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[9]~1 (
	.dataa(state_4),
	.datab(\count[8]~q ),
	.datac(\state~q ),
	.datad(\count[9]~0_combout ),
	.cin(gnd),
	.combout(\count[9]~1_combout ),
	.cout());
defparam \count[9]~1 .lut_mask = 16'hF7FF;
defparam \count[9]~1 .sum_lutc_input = "datac";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cycloneive_lcell_comb \count~4 (
	.dataa(state_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hAAFF;
defparam \count~4 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \wdata[1]~0 (
	.dataa(\state~q ),
	.datab(state_4),
	.datac(splitter_nodes_receive_0_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\wdata[1]~0_combout ),
	.cout());
defparam \wdata[1]~0 .lut_mask = 16'hFEFF;
defparam \wdata[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \user_saw_rvalid~0 (
	.dataa(\td_shift[0]~q ),
	.datab(\user_saw_rvalid~q ),
	.datac(irf_reg_0_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.cout());
defparam \user_saw_rvalid~0 .lut_mask = 16'hACAC;
defparam \user_saw_rvalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \user_saw_rvalid~1 (
	.dataa(\user_saw_rvalid~q ),
	.datab(\count[0]~q ),
	.datac(\wdata[1]~0_combout ),
	.datad(\user_saw_rvalid~0_combout ),
	.cin(gnd),
	.combout(\user_saw_rvalid~1_combout ),
	.cout());
defparam \user_saw_rvalid~1 .lut_mask = 16'hFFBE;
defparam \user_saw_rvalid~1 .sum_lutc_input = "datac";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~11 (
	.dataa(altera_internal_jtag1),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~11_combout ),
	.cout());
defparam \td_shift~11 .lut_mask = 16'hEEEE;
defparam \td_shift~11 .sum_lutc_input = "datac";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cycloneive_lcell_comb \r_ena~0 (
	.dataa(r_val),
	.datab(r_ena11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\r_ena~0_combout ),
	.cout());
defparam \r_ena~0 .lut_mask = 16'hEEEE;
defparam \r_ena~0 .sum_lutc_input = "datac";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cycloneive_lcell_comb \td_shift~8 (
	.dataa(\td_shift[10]~q ),
	.datab(\rdata[7]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~8_combout ),
	.cout());
defparam \td_shift~8 .lut_mask = 16'hAACC;
defparam \td_shift~8 .sum_lutc_input = "datac";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cycloneive_lcell_comb \td_shift~6 (
	.dataa(\user_saw_rvalid~q ),
	.datab(\td_shift[9]~q ),
	.datac(\state~q ),
	.datad(\count[1]~q ),
	.cin(gnd),
	.combout(\td_shift~6_combout ),
	.cout());
defparam \td_shift~6 .lut_mask = 16'hEFFF;
defparam \td_shift~6 .sum_lutc_input = "datac";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cycloneive_lcell_comb \td_shift~22 (
	.dataa(\td_shift[9]~q ),
	.datab(\rdata[6]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~22_combout ),
	.cout());
defparam \td_shift~22 .lut_mask = 16'hAACC;
defparam \td_shift~22 .sum_lutc_input = "datac";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~22_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cycloneive_lcell_comb \td_shift~20 (
	.dataa(\td_shift[8]~q ),
	.datab(\rdata[5]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~20_combout ),
	.cout());
defparam \td_shift~20 .lut_mask = 16'hACAC;
defparam \td_shift~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~21 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(\td_shift~20_combout ),
	.cin(gnd),
	.combout(\td_shift~21_combout ),
	.cout());
defparam \td_shift~21 .lut_mask = 16'hFFFE;
defparam \td_shift~21 .sum_lutc_input = "datac";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~21_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cycloneive_lcell_comb \td_shift~18 (
	.dataa(\td_shift[7]~q ),
	.datab(\rdata[4]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~18_combout ),
	.cout());
defparam \td_shift~18 .lut_mask = 16'hAACC;
defparam \td_shift~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~19 (
	.dataa(\td_shift~18_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~19_combout ),
	.cout());
defparam \td_shift~19 .lut_mask = 16'hFAFC;
defparam \td_shift~19 .sum_lutc_input = "datac";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~19_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cycloneive_lcell_comb \td_shift~16 (
	.dataa(\td_shift[6]~q ),
	.datab(\rdata[3]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~16_combout ),
	.cout());
defparam \td_shift~16 .lut_mask = 16'hAACC;
defparam \td_shift~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~17 (
	.dataa(\td_shift~16_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~17_combout ),
	.cout());
defparam \td_shift~17 .lut_mask = 16'hFAFC;
defparam \td_shift~17 .sum_lutc_input = "datac";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~17_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cycloneive_lcell_comb \td_shift~14 (
	.dataa(\td_shift[5]~q ),
	.datab(\rdata[2]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~14_combout ),
	.cout());
defparam \td_shift~14 .lut_mask = 16'hACAC;
defparam \td_shift~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~15 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(\td_shift~14_combout ),
	.cin(gnd),
	.combout(\td_shift~15_combout ),
	.cout());
defparam \td_shift~15 .lut_mask = 16'hFFFE;
defparam \td_shift~15 .sum_lutc_input = "datac";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~15_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cycloneive_lcell_comb \td_shift~12 (
	.dataa(\td_shift[4]~q ),
	.datab(\rdata[1]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~12_combout ),
	.cout());
defparam \td_shift~12 .lut_mask = 16'hACAC;
defparam \td_shift~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~13 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(\td_shift~12_combout ),
	.cin(gnd),
	.combout(\td_shift~13_combout ),
	.cout());
defparam \td_shift~13 .lut_mask = 16'hFFFE;
defparam \td_shift~13 .sum_lutc_input = "datac";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~13_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

cycloneive_lcell_comb \td_shift~9 (
	.dataa(\td_shift[3]~q ),
	.datab(\rdata[0]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~9_combout ),
	.cout());
defparam \td_shift~9 .lut_mask = 16'hAACC;
defparam \td_shift~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~10 (
	.dataa(\td_shift~9_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~10_combout ),
	.cout());
defparam \td_shift~10 .lut_mask = 16'hFAFC;
defparam \td_shift~10 .sum_lutc_input = "datac";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cycloneive_lcell_comb \write_stalled~0 (
	.dataa(\td_shift[10]~q ),
	.datab(\write_stalled~q ),
	.datac(\tck_t_dav~q ),
	.datad(altera_internal_jtag1),
	.cin(gnd),
	.combout(\write_stalled~0_combout ),
	.cout());
defparam \write_stalled~0 .lut_mask = 16'hEFFF;
defparam \write_stalled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~1 (
	.dataa(state_4),
	.datab(splitter_nodes_receive_0_3),
	.datac(virtual_ir_scan_reg),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_stalled~1_combout ),
	.cout());
defparam \write_stalled~1 .lut_mask = 16'hEFEF;
defparam \write_stalled~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~2 (
	.dataa(\count[1]~q ),
	.datab(irf_reg_0_1),
	.datac(\state~q ),
	.datad(\write_stalled~1_combout ),
	.cin(gnd),
	.combout(\write_stalled~2_combout ),
	.cout());
defparam \write_stalled~2 .lut_mask = 16'hFFFB;
defparam \write_stalled~2 .sum_lutc_input = "datac";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cycloneive_lcell_comb \td_shift~5 (
	.dataa(\td_shift[2]~q ),
	.datab(\write_stalled~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~5_combout ),
	.cout());
defparam \td_shift~5 .lut_mask = 16'hAACC;
defparam \td_shift~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~7 (
	.dataa(\td_shift~5_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~7_combout ),
	.cout());
defparam \td_shift~7 .lut_mask = 16'hFAFC;
defparam \td_shift~7 .sum_lutc_input = "datac";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~0 (
	.dataa(\td_shift[1]~q ),
	.datab(\rvalid~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~0_combout ),
	.cout());
defparam \td_shift~0 .lut_mask = 16'hACAC;
defparam \td_shift~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~1 (
	.dataa(\user_saw_rvalid~q ),
	.datab(\td_shift[9]~q ),
	.datac(\count[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~1_combout ),
	.cout());
defparam \td_shift~1 .lut_mask = 16'hF7F7;
defparam \td_shift~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~2 (
	.dataa(\state~q ),
	.datab(altera_internal_jtag1),
	.datac(irf_reg_0_1),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~2_combout ),
	.cout());
defparam \td_shift~2 .lut_mask = 16'hDF8F;
defparam \td_shift~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~3 (
	.dataa(\tck_t_dav~q ),
	.datab(\td_shift~0_combout ),
	.datac(\state~q ),
	.datad(\td_shift~2_combout ),
	.cin(gnd),
	.combout(\td_shift~3_combout ),
	.cout());
defparam \td_shift~3 .lut_mask = 16'hAFCF;
defparam \td_shift~3 .sum_lutc_input = "datac";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cycloneive_lcell_comb \rvalid0~0 (
	.dataa(rvalid01),
	.datab(r_val),
	.datac(r_ena11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rvalid0~0_combout ),
	.cout());
defparam \rvalid0~0 .lut_mask = 16'h7F7F;
defparam \rvalid0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h5555;
defparam \read~0 .sum_lutc_input = "datac";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cycloneive_lcell_comb \rvalid0~1 (
	.dataa(\read1~q ),
	.datab(\read2~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\read_req~q ),
	.cin(gnd),
	.combout(\rvalid0~1_combout ),
	.cout());
defparam \rvalid0~1 .lut_mask = 16'h6FFF;
defparam \rvalid0~1 .sum_lutc_input = "datac";

dffeas rst2(
	.clk(clk),
	.d(sink_in_reset),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cycloneive_lcell_comb \rvalid0~2 (
	.dataa(\rvalid0~0_combout ),
	.datab(\rvalid0~1_combout ),
	.datac(gnd),
	.datad(\rst2~q ),
	.cin(gnd),
	.combout(\rvalid0~2_combout ),
	.cout());
defparam \rvalid0~2 .lut_mask = 16'hDDFF;
defparam \rvalid0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~0 (
	.dataa(\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'h5555;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wdata[1]~1 (
	.dataa(\count[8]~q ),
	.datab(irf_reg_0_1),
	.datac(\state~q ),
	.datad(\write_stalled~1_combout ),
	.cin(gnd),
	.combout(\wdata[1]~1_combout ),
	.cout());
defparam \wdata[1]~1 .lut_mask = 16'hFFFB;
defparam \wdata[1]~1 .sum_lutc_input = "datac";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cycloneive_lcell_comb \always2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\write1~q ),
	.datad(\write2~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h0FF0;
defparam \always2~0 .sum_lutc_input = "datac";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cycloneive_lcell_comb \t_pause~0 (
	.dataa(\always2~0_combout ),
	.datab(t_dav),
	.datac(\write_stalled~q ),
	.datad(\write_valid~q ),
	.cin(gnd),
	.combout(\t_pause~0_combout ),
	.cout());
defparam \t_pause~0 .lut_mask = 16'hFEFF;
defparam \t_pause~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jupdate~0 (
	.dataa(\jupdate~q ),
	.datab(irf_reg_0_1),
	.datac(\always0~0_combout ),
	.datad(state_8),
	.cin(gnd),
	.combout(\jupdate~0_combout ),
	.cout());
defparam \jupdate~0 .lut_mask = 16'h6996;
defparam \jupdate~0 .sum_lutc_input = "datac";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cycloneive_lcell_comb \t_pause~1 (
	.dataa(\rst2~q ),
	.datab(\t_pause~0_combout ),
	.datac(\jupdate1~q ),
	.datad(\jupdate2~q ),
	.cin(gnd),
	.combout(\t_pause~1_combout ),
	.cout());
defparam \t_pause~1 .lut_mask = 16'hEFFE;
defparam \t_pause~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_ena~2 (
	.dataa(t_ena1),
	.datab(\write_valid~q ),
	.datac(t_dav),
	.datad(\write_stalled~q ),
	.cin(gnd),
	.combout(\t_ena~2_combout ),
	.cout());
defparam \t_ena~2 .lut_mask = 16'hEFFF;
defparam \t_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_ena~3 (
	.dataa(\write1~q ),
	.datab(\write2~q ),
	.datac(\rst2~q ),
	.datad(\t_ena~2_combout ),
	.cin(gnd),
	.combout(\t_ena~3_combout ),
	.cout());
defparam \t_ena~3 .lut_mask = 16'hFFF6;
defparam \t_ena~3 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_jtag_uart_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	rvalid,
	wr_rfifo,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	rvalid;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_6;
input 	wdata_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.rvalid(rvalid),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module usb_system_scfifo_1 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	rvalid,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	rvalid;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_scfifo_jr21 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.rvalid(rvalid),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module usb_system_scfifo_jr21 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	rvalid,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	rvalid;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_a_dpfifo_q131 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.rvalid(rvalid),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module usb_system_a_dpfifo_q131 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	rvalid,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	rvalid;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


usb_system_cntr_1ob_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

usb_system_cntr_1ob rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.rvalid(rvalid),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

usb_system_dpram_nl21 FIFOram(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.outclocken(rvalid),
	.wren(wreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wraddress({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.rdaddress({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.outclock(clock));

usb_system_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.rvalid(rvalid),
	.wreq(wreq),
	.clock(clock));

endmodule

module usb_system_a_fefifo_7cf (
	r_sync_rst,
	b_full1,
	b_non_empty1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	rvalid,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	b_non_empty1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	rvalid;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \b_non_empty~1_combout ;


usb_system_cntr_do7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.updown(wreq),
	._(\_~4_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~4 (
	.dataa(t_ena),
	.datab(b_full1),
	.datac(rvalid),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'h9696;
defparam \_~4 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cycloneive_lcell_comb \b_full~0 (
	.dataa(b_non_empty1),
	.datab(counter_reg_bit_3),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_1),
	.datad(t_ena),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(rvalid),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(b_full1),
	.datab(t_ena),
	.datac(gnd),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hEEFF;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_4),
	.datab(counter_reg_bit_5),
	.datac(wreq),
	.datad(\_~2_combout ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFFFE;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(\b_non_empty~0_combout ),
	.datab(b_non_empty1),
	.datac(\_~3_combout ),
	.datad(rvalid),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hFEFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

endmodule

module usb_system_cntr_do7 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module usb_system_cntr_1ob (
	r_sync_rst,
	rvalid,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	rvalid;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rvalid),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module usb_system_cntr_1ob_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module usb_system_dpram_nl21 (
	q,
	outclocken,
	wren,
	data,
	wraddress,
	rdaddress,
	outclock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	outclocken;
input 	wren;
input 	[7:0] data;
input 	[5:0] wraddress;
input 	[5:0] rdaddress;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_r1m1 altsyncram1(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(outclocken),
	.wren_a(wren),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({wraddress[5],wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.address_b({rdaddress[5],rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.clock1(outclock),
	.clock0(outclock));

endmodule

module usb_system_altsyncram_r1m1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block2a0_PORTBDATAOUT_bus;
wire [143:0] ram_block2a1_PORTBDATAOUT_bus;
wire [143:0] ram_block2a2_PORTBDATAOUT_bus;
wire [143:0] ram_block2a3_PORTBDATAOUT_bus;
wire [143:0] ram_block2a4_PORTBDATAOUT_bus;
wire [143:0] ram_block2a5_PORTBDATAOUT_bus;
wire [143:0] ram_block2a6_PORTBDATAOUT_bus;
wire [143:0] ram_block2a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block2a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block2a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block2a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block2a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block2a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block2a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block2a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block2a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block2a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a0_PORTBDATAOUT_bus));
defparam ram_block2a0.clk0_core_clock_enable = "ena0";
defparam ram_block2a0.clk1_core_clock_enable = "ena1";
defparam ram_block2a0.clk1_input_clock_enable = "ena1";
defparam ram_block2a0.data_interleave_offset_in_bits = 1;
defparam ram_block2a0.data_interleave_width_in_bits = 1;
defparam ram_block2a0.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a0.operation_mode = "dual_port";
defparam ram_block2a0.port_a_address_clear = "none";
defparam ram_block2a0.port_a_address_width = 6;
defparam ram_block2a0.port_a_data_out_clear = "none";
defparam ram_block2a0.port_a_data_out_clock = "none";
defparam ram_block2a0.port_a_data_width = 1;
defparam ram_block2a0.port_a_first_address = 0;
defparam ram_block2a0.port_a_first_bit_number = 0;
defparam ram_block2a0.port_a_last_address = 63;
defparam ram_block2a0.port_a_logical_ram_depth = 64;
defparam ram_block2a0.port_a_logical_ram_width = 8;
defparam ram_block2a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_address_clear = "none";
defparam ram_block2a0.port_b_address_clock = "clock1";
defparam ram_block2a0.port_b_address_width = 6;
defparam ram_block2a0.port_b_data_out_clear = "none";
defparam ram_block2a0.port_b_data_out_clock = "none";
defparam ram_block2a0.port_b_data_width = 1;
defparam ram_block2a0.port_b_first_address = 0;
defparam ram_block2a0.port_b_first_bit_number = 0;
defparam ram_block2a0.port_b_last_address = 63;
defparam ram_block2a0.port_b_logical_ram_depth = 64;
defparam ram_block2a0.port_b_logical_ram_width = 8;
defparam ram_block2a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_read_enable_clock = "clock1";
defparam ram_block2a0.ram_block_type = "auto";

cycloneive_ram_block ram_block2a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a1_PORTBDATAOUT_bus));
defparam ram_block2a1.clk0_core_clock_enable = "ena0";
defparam ram_block2a1.clk1_core_clock_enable = "ena1";
defparam ram_block2a1.clk1_input_clock_enable = "ena1";
defparam ram_block2a1.data_interleave_offset_in_bits = 1;
defparam ram_block2a1.data_interleave_width_in_bits = 1;
defparam ram_block2a1.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a1.operation_mode = "dual_port";
defparam ram_block2a1.port_a_address_clear = "none";
defparam ram_block2a1.port_a_address_width = 6;
defparam ram_block2a1.port_a_data_out_clear = "none";
defparam ram_block2a1.port_a_data_out_clock = "none";
defparam ram_block2a1.port_a_data_width = 1;
defparam ram_block2a1.port_a_first_address = 0;
defparam ram_block2a1.port_a_first_bit_number = 1;
defparam ram_block2a1.port_a_last_address = 63;
defparam ram_block2a1.port_a_logical_ram_depth = 64;
defparam ram_block2a1.port_a_logical_ram_width = 8;
defparam ram_block2a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_address_clear = "none";
defparam ram_block2a1.port_b_address_clock = "clock1";
defparam ram_block2a1.port_b_address_width = 6;
defparam ram_block2a1.port_b_data_out_clear = "none";
defparam ram_block2a1.port_b_data_out_clock = "none";
defparam ram_block2a1.port_b_data_width = 1;
defparam ram_block2a1.port_b_first_address = 0;
defparam ram_block2a1.port_b_first_bit_number = 1;
defparam ram_block2a1.port_b_last_address = 63;
defparam ram_block2a1.port_b_logical_ram_depth = 64;
defparam ram_block2a1.port_b_logical_ram_width = 8;
defparam ram_block2a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_read_enable_clock = "clock1";
defparam ram_block2a1.ram_block_type = "auto";

cycloneive_ram_block ram_block2a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a2_PORTBDATAOUT_bus));
defparam ram_block2a2.clk0_core_clock_enable = "ena0";
defparam ram_block2a2.clk1_core_clock_enable = "ena1";
defparam ram_block2a2.clk1_input_clock_enable = "ena1";
defparam ram_block2a2.data_interleave_offset_in_bits = 1;
defparam ram_block2a2.data_interleave_width_in_bits = 1;
defparam ram_block2a2.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a2.operation_mode = "dual_port";
defparam ram_block2a2.port_a_address_clear = "none";
defparam ram_block2a2.port_a_address_width = 6;
defparam ram_block2a2.port_a_data_out_clear = "none";
defparam ram_block2a2.port_a_data_out_clock = "none";
defparam ram_block2a2.port_a_data_width = 1;
defparam ram_block2a2.port_a_first_address = 0;
defparam ram_block2a2.port_a_first_bit_number = 2;
defparam ram_block2a2.port_a_last_address = 63;
defparam ram_block2a2.port_a_logical_ram_depth = 64;
defparam ram_block2a2.port_a_logical_ram_width = 8;
defparam ram_block2a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_address_clear = "none";
defparam ram_block2a2.port_b_address_clock = "clock1";
defparam ram_block2a2.port_b_address_width = 6;
defparam ram_block2a2.port_b_data_out_clear = "none";
defparam ram_block2a2.port_b_data_out_clock = "none";
defparam ram_block2a2.port_b_data_width = 1;
defparam ram_block2a2.port_b_first_address = 0;
defparam ram_block2a2.port_b_first_bit_number = 2;
defparam ram_block2a2.port_b_last_address = 63;
defparam ram_block2a2.port_b_logical_ram_depth = 64;
defparam ram_block2a2.port_b_logical_ram_width = 8;
defparam ram_block2a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_read_enable_clock = "clock1";
defparam ram_block2a2.ram_block_type = "auto";

cycloneive_ram_block ram_block2a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a3_PORTBDATAOUT_bus));
defparam ram_block2a3.clk0_core_clock_enable = "ena0";
defparam ram_block2a3.clk1_core_clock_enable = "ena1";
defparam ram_block2a3.clk1_input_clock_enable = "ena1";
defparam ram_block2a3.data_interleave_offset_in_bits = 1;
defparam ram_block2a3.data_interleave_width_in_bits = 1;
defparam ram_block2a3.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a3.operation_mode = "dual_port";
defparam ram_block2a3.port_a_address_clear = "none";
defparam ram_block2a3.port_a_address_width = 6;
defparam ram_block2a3.port_a_data_out_clear = "none";
defparam ram_block2a3.port_a_data_out_clock = "none";
defparam ram_block2a3.port_a_data_width = 1;
defparam ram_block2a3.port_a_first_address = 0;
defparam ram_block2a3.port_a_first_bit_number = 3;
defparam ram_block2a3.port_a_last_address = 63;
defparam ram_block2a3.port_a_logical_ram_depth = 64;
defparam ram_block2a3.port_a_logical_ram_width = 8;
defparam ram_block2a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_address_clear = "none";
defparam ram_block2a3.port_b_address_clock = "clock1";
defparam ram_block2a3.port_b_address_width = 6;
defparam ram_block2a3.port_b_data_out_clear = "none";
defparam ram_block2a3.port_b_data_out_clock = "none";
defparam ram_block2a3.port_b_data_width = 1;
defparam ram_block2a3.port_b_first_address = 0;
defparam ram_block2a3.port_b_first_bit_number = 3;
defparam ram_block2a3.port_b_last_address = 63;
defparam ram_block2a3.port_b_logical_ram_depth = 64;
defparam ram_block2a3.port_b_logical_ram_width = 8;
defparam ram_block2a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_read_enable_clock = "clock1";
defparam ram_block2a3.ram_block_type = "auto";

cycloneive_ram_block ram_block2a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a4_PORTBDATAOUT_bus));
defparam ram_block2a4.clk0_core_clock_enable = "ena0";
defparam ram_block2a4.clk1_core_clock_enable = "ena1";
defparam ram_block2a4.clk1_input_clock_enable = "ena1";
defparam ram_block2a4.data_interleave_offset_in_bits = 1;
defparam ram_block2a4.data_interleave_width_in_bits = 1;
defparam ram_block2a4.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a4.operation_mode = "dual_port";
defparam ram_block2a4.port_a_address_clear = "none";
defparam ram_block2a4.port_a_address_width = 6;
defparam ram_block2a4.port_a_data_out_clear = "none";
defparam ram_block2a4.port_a_data_out_clock = "none";
defparam ram_block2a4.port_a_data_width = 1;
defparam ram_block2a4.port_a_first_address = 0;
defparam ram_block2a4.port_a_first_bit_number = 4;
defparam ram_block2a4.port_a_last_address = 63;
defparam ram_block2a4.port_a_logical_ram_depth = 64;
defparam ram_block2a4.port_a_logical_ram_width = 8;
defparam ram_block2a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_address_clear = "none";
defparam ram_block2a4.port_b_address_clock = "clock1";
defparam ram_block2a4.port_b_address_width = 6;
defparam ram_block2a4.port_b_data_out_clear = "none";
defparam ram_block2a4.port_b_data_out_clock = "none";
defparam ram_block2a4.port_b_data_width = 1;
defparam ram_block2a4.port_b_first_address = 0;
defparam ram_block2a4.port_b_first_bit_number = 4;
defparam ram_block2a4.port_b_last_address = 63;
defparam ram_block2a4.port_b_logical_ram_depth = 64;
defparam ram_block2a4.port_b_logical_ram_width = 8;
defparam ram_block2a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_read_enable_clock = "clock1";
defparam ram_block2a4.ram_block_type = "auto";

cycloneive_ram_block ram_block2a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a5_PORTBDATAOUT_bus));
defparam ram_block2a5.clk0_core_clock_enable = "ena0";
defparam ram_block2a5.clk1_core_clock_enable = "ena1";
defparam ram_block2a5.clk1_input_clock_enable = "ena1";
defparam ram_block2a5.data_interleave_offset_in_bits = 1;
defparam ram_block2a5.data_interleave_width_in_bits = 1;
defparam ram_block2a5.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a5.operation_mode = "dual_port";
defparam ram_block2a5.port_a_address_clear = "none";
defparam ram_block2a5.port_a_address_width = 6;
defparam ram_block2a5.port_a_data_out_clear = "none";
defparam ram_block2a5.port_a_data_out_clock = "none";
defparam ram_block2a5.port_a_data_width = 1;
defparam ram_block2a5.port_a_first_address = 0;
defparam ram_block2a5.port_a_first_bit_number = 5;
defparam ram_block2a5.port_a_last_address = 63;
defparam ram_block2a5.port_a_logical_ram_depth = 64;
defparam ram_block2a5.port_a_logical_ram_width = 8;
defparam ram_block2a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_address_clear = "none";
defparam ram_block2a5.port_b_address_clock = "clock1";
defparam ram_block2a5.port_b_address_width = 6;
defparam ram_block2a5.port_b_data_out_clear = "none";
defparam ram_block2a5.port_b_data_out_clock = "none";
defparam ram_block2a5.port_b_data_width = 1;
defparam ram_block2a5.port_b_first_address = 0;
defparam ram_block2a5.port_b_first_bit_number = 5;
defparam ram_block2a5.port_b_last_address = 63;
defparam ram_block2a5.port_b_logical_ram_depth = 64;
defparam ram_block2a5.port_b_logical_ram_width = 8;
defparam ram_block2a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_read_enable_clock = "clock1";
defparam ram_block2a5.ram_block_type = "auto";

cycloneive_ram_block ram_block2a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a6_PORTBDATAOUT_bus));
defparam ram_block2a6.clk0_core_clock_enable = "ena0";
defparam ram_block2a6.clk1_core_clock_enable = "ena1";
defparam ram_block2a6.clk1_input_clock_enable = "ena1";
defparam ram_block2a6.data_interleave_offset_in_bits = 1;
defparam ram_block2a6.data_interleave_width_in_bits = 1;
defparam ram_block2a6.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a6.operation_mode = "dual_port";
defparam ram_block2a6.port_a_address_clear = "none";
defparam ram_block2a6.port_a_address_width = 6;
defparam ram_block2a6.port_a_data_out_clear = "none";
defparam ram_block2a6.port_a_data_out_clock = "none";
defparam ram_block2a6.port_a_data_width = 1;
defparam ram_block2a6.port_a_first_address = 0;
defparam ram_block2a6.port_a_first_bit_number = 6;
defparam ram_block2a6.port_a_last_address = 63;
defparam ram_block2a6.port_a_logical_ram_depth = 64;
defparam ram_block2a6.port_a_logical_ram_width = 8;
defparam ram_block2a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_address_clear = "none";
defparam ram_block2a6.port_b_address_clock = "clock1";
defparam ram_block2a6.port_b_address_width = 6;
defparam ram_block2a6.port_b_data_out_clear = "none";
defparam ram_block2a6.port_b_data_out_clock = "none";
defparam ram_block2a6.port_b_data_width = 1;
defparam ram_block2a6.port_b_first_address = 0;
defparam ram_block2a6.port_b_first_bit_number = 6;
defparam ram_block2a6.port_b_last_address = 63;
defparam ram_block2a6.port_b_logical_ram_depth = 64;
defparam ram_block2a6.port_b_logical_ram_width = 8;
defparam ram_block2a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_read_enable_clock = "clock1";
defparam ram_block2a6.ram_block_type = "auto";

cycloneive_ram_block ram_block2a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a7_PORTBDATAOUT_bus));
defparam ram_block2a7.clk0_core_clock_enable = "ena0";
defparam ram_block2a7.clk1_core_clock_enable = "ena1";
defparam ram_block2a7.clk1_input_clock_enable = "ena1";
defparam ram_block2a7.data_interleave_offset_in_bits = 1;
defparam ram_block2a7.data_interleave_width_in_bits = 1;
defparam ram_block2a7.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_r:the_usb_system_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a7.operation_mode = "dual_port";
defparam ram_block2a7.port_a_address_clear = "none";
defparam ram_block2a7.port_a_address_width = 6;
defparam ram_block2a7.port_a_data_out_clear = "none";
defparam ram_block2a7.port_a_data_out_clock = "none";
defparam ram_block2a7.port_a_data_width = 1;
defparam ram_block2a7.port_a_first_address = 0;
defparam ram_block2a7.port_a_first_bit_number = 7;
defparam ram_block2a7.port_a_last_address = 63;
defparam ram_block2a7.port_a_logical_ram_depth = 64;
defparam ram_block2a7.port_a_logical_ram_width = 8;
defparam ram_block2a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_address_clear = "none";
defparam ram_block2a7.port_b_address_clock = "clock1";
defparam ram_block2a7.port_b_address_width = 6;
defparam ram_block2a7.port_b_data_out_clear = "none";
defparam ram_block2a7.port_b_data_out_clock = "none";
defparam ram_block2a7.port_b_data_width = 1;
defparam ram_block2a7.port_b_first_address = 0;
defparam ram_block2a7.port_b_first_bit_number = 7;
defparam ram_block2a7.port_b_last_address = 63;
defparam ram_block2a7.port_b_logical_ram_depth = 64;
defparam ram_block2a7.port_b_logical_ram_width = 8;
defparam ram_block2a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_read_enable_clock = "clock1";
defparam ram_block2a7.ram_block_type = "auto";

endmodule

module usb_system_usb_system_jtag_uart_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	fifo_wr,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	fifo_wr;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(fifo_wr),
	.clock(clk_clk));

endmodule

module usb_system_scfifo_2 (
	q,
	data,
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	wrreq,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_scfifo_jr21_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(wrreq),
	.clock(clock));

endmodule

module usb_system_scfifo_jr21_1 (
	q,
	data,
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	wrreq,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_a_dpfifo_q131_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wreq(wrreq),
	.clock(clock));

endmodule

module usb_system_a_dpfifo_q131_1 (
	q,
	data,
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


usb_system_cntr_1ob_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

usb_system_cntr_1ob_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

usb_system_dpram_nl21_1 FIFOram(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.outclocken(r_val),
	.wren(wreq),
	.wraddress({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.rdaddress({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.outclock(clock));

usb_system_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full1(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.wreq(wreq),
	.clock(clock));

endmodule

module usb_system_a_fefifo_7cf_1 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty1,
	r_val,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty1;
input 	r_val;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;


usb_system_cntr_do7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.updown(wreq),
	._(\_~0_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(wreq),
	.datad(r_val),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FF0;
defparam \_~0 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cycloneive_lcell_comb \b_full~0 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(wreq),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hFFFE;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(counter_reg_bit_3),
	.datab(\b_non_empty~0_combout ),
	.datac(counter_reg_bit_0),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hEFFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~2 (
	.dataa(b_full1),
	.datab(wreq),
	.datac(b_non_empty1),
	.datad(\b_non_empty~1_combout ),
	.cin(gnd),
	.combout(\b_non_empty~2_combout ),
	.cout());
defparam \b_non_empty~2 .lut_mask = 16'hFFFE;
defparam \b_non_empty~2 .sum_lutc_input = "datac";

endmodule

module usb_system_cntr_do7_1 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module usb_system_cntr_1ob_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module usb_system_cntr_1ob_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module usb_system_dpram_nl21_1 (
	q,
	data,
	outclocken,
	wren,
	wraddress,
	rdaddress,
	outclock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	outclocken;
input 	wren;
input 	[5:0] wraddress;
input 	[5:0] rdaddress;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altsyncram_r1m1_1 altsyncram1(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clocken1(outclocken),
	.wren_a(wren),
	.address_a({wraddress[5],wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.address_b({rdaddress[5],rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.clock1(outclock),
	.clock0(outclock));

endmodule

module usb_system_altsyncram_r1m1_1 (
	q_b,
	data_a,
	clocken1,
	wren_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	clocken1;
input 	wren_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block2a7_PORTBDATAOUT_bus;
wire [143:0] ram_block2a0_PORTBDATAOUT_bus;
wire [143:0] ram_block2a1_PORTBDATAOUT_bus;
wire [143:0] ram_block2a2_PORTBDATAOUT_bus;
wire [143:0] ram_block2a3_PORTBDATAOUT_bus;
wire [143:0] ram_block2a4_PORTBDATAOUT_bus;
wire [143:0] ram_block2a5_PORTBDATAOUT_bus;
wire [143:0] ram_block2a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block2a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block2a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block2a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block2a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block2a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block2a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block2a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block2a6_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block2a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a7_PORTBDATAOUT_bus));
defparam ram_block2a7.clk0_core_clock_enable = "ena0";
defparam ram_block2a7.clk1_core_clock_enable = "ena1";
defparam ram_block2a7.clk1_input_clock_enable = "ena1";
defparam ram_block2a7.data_interleave_offset_in_bits = 1;
defparam ram_block2a7.data_interleave_width_in_bits = 1;
defparam ram_block2a7.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a7.operation_mode = "dual_port";
defparam ram_block2a7.port_a_address_clear = "none";
defparam ram_block2a7.port_a_address_width = 6;
defparam ram_block2a7.port_a_data_out_clear = "none";
defparam ram_block2a7.port_a_data_out_clock = "none";
defparam ram_block2a7.port_a_data_width = 1;
defparam ram_block2a7.port_a_first_address = 0;
defparam ram_block2a7.port_a_first_bit_number = 7;
defparam ram_block2a7.port_a_last_address = 63;
defparam ram_block2a7.port_a_logical_ram_depth = 64;
defparam ram_block2a7.port_a_logical_ram_width = 8;
defparam ram_block2a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_address_clear = "none";
defparam ram_block2a7.port_b_address_clock = "clock1";
defparam ram_block2a7.port_b_address_width = 6;
defparam ram_block2a7.port_b_data_out_clear = "none";
defparam ram_block2a7.port_b_data_out_clock = "none";
defparam ram_block2a7.port_b_data_width = 1;
defparam ram_block2a7.port_b_first_address = 0;
defparam ram_block2a7.port_b_first_bit_number = 7;
defparam ram_block2a7.port_b_last_address = 63;
defparam ram_block2a7.port_b_logical_ram_depth = 64;
defparam ram_block2a7.port_b_logical_ram_width = 8;
defparam ram_block2a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_read_enable_clock = "clock1";
defparam ram_block2a7.ram_block_type = "auto";

cycloneive_ram_block ram_block2a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a0_PORTBDATAOUT_bus));
defparam ram_block2a0.clk0_core_clock_enable = "ena0";
defparam ram_block2a0.clk1_core_clock_enable = "ena1";
defparam ram_block2a0.clk1_input_clock_enable = "ena1";
defparam ram_block2a0.data_interleave_offset_in_bits = 1;
defparam ram_block2a0.data_interleave_width_in_bits = 1;
defparam ram_block2a0.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a0.operation_mode = "dual_port";
defparam ram_block2a0.port_a_address_clear = "none";
defparam ram_block2a0.port_a_address_width = 6;
defparam ram_block2a0.port_a_data_out_clear = "none";
defparam ram_block2a0.port_a_data_out_clock = "none";
defparam ram_block2a0.port_a_data_width = 1;
defparam ram_block2a0.port_a_first_address = 0;
defparam ram_block2a0.port_a_first_bit_number = 0;
defparam ram_block2a0.port_a_last_address = 63;
defparam ram_block2a0.port_a_logical_ram_depth = 64;
defparam ram_block2a0.port_a_logical_ram_width = 8;
defparam ram_block2a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_address_clear = "none";
defparam ram_block2a0.port_b_address_clock = "clock1";
defparam ram_block2a0.port_b_address_width = 6;
defparam ram_block2a0.port_b_data_out_clear = "none";
defparam ram_block2a0.port_b_data_out_clock = "none";
defparam ram_block2a0.port_b_data_width = 1;
defparam ram_block2a0.port_b_first_address = 0;
defparam ram_block2a0.port_b_first_bit_number = 0;
defparam ram_block2a0.port_b_last_address = 63;
defparam ram_block2a0.port_b_logical_ram_depth = 64;
defparam ram_block2a0.port_b_logical_ram_width = 8;
defparam ram_block2a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_read_enable_clock = "clock1";
defparam ram_block2a0.ram_block_type = "auto";

cycloneive_ram_block ram_block2a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a1_PORTBDATAOUT_bus));
defparam ram_block2a1.clk0_core_clock_enable = "ena0";
defparam ram_block2a1.clk1_core_clock_enable = "ena1";
defparam ram_block2a1.clk1_input_clock_enable = "ena1";
defparam ram_block2a1.data_interleave_offset_in_bits = 1;
defparam ram_block2a1.data_interleave_width_in_bits = 1;
defparam ram_block2a1.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a1.operation_mode = "dual_port";
defparam ram_block2a1.port_a_address_clear = "none";
defparam ram_block2a1.port_a_address_width = 6;
defparam ram_block2a1.port_a_data_out_clear = "none";
defparam ram_block2a1.port_a_data_out_clock = "none";
defparam ram_block2a1.port_a_data_width = 1;
defparam ram_block2a1.port_a_first_address = 0;
defparam ram_block2a1.port_a_first_bit_number = 1;
defparam ram_block2a1.port_a_last_address = 63;
defparam ram_block2a1.port_a_logical_ram_depth = 64;
defparam ram_block2a1.port_a_logical_ram_width = 8;
defparam ram_block2a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_address_clear = "none";
defparam ram_block2a1.port_b_address_clock = "clock1";
defparam ram_block2a1.port_b_address_width = 6;
defparam ram_block2a1.port_b_data_out_clear = "none";
defparam ram_block2a1.port_b_data_out_clock = "none";
defparam ram_block2a1.port_b_data_width = 1;
defparam ram_block2a1.port_b_first_address = 0;
defparam ram_block2a1.port_b_first_bit_number = 1;
defparam ram_block2a1.port_b_last_address = 63;
defparam ram_block2a1.port_b_logical_ram_depth = 64;
defparam ram_block2a1.port_b_logical_ram_width = 8;
defparam ram_block2a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_read_enable_clock = "clock1";
defparam ram_block2a1.ram_block_type = "auto";

cycloneive_ram_block ram_block2a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a2_PORTBDATAOUT_bus));
defparam ram_block2a2.clk0_core_clock_enable = "ena0";
defparam ram_block2a2.clk1_core_clock_enable = "ena1";
defparam ram_block2a2.clk1_input_clock_enable = "ena1";
defparam ram_block2a2.data_interleave_offset_in_bits = 1;
defparam ram_block2a2.data_interleave_width_in_bits = 1;
defparam ram_block2a2.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a2.operation_mode = "dual_port";
defparam ram_block2a2.port_a_address_clear = "none";
defparam ram_block2a2.port_a_address_width = 6;
defparam ram_block2a2.port_a_data_out_clear = "none";
defparam ram_block2a2.port_a_data_out_clock = "none";
defparam ram_block2a2.port_a_data_width = 1;
defparam ram_block2a2.port_a_first_address = 0;
defparam ram_block2a2.port_a_first_bit_number = 2;
defparam ram_block2a2.port_a_last_address = 63;
defparam ram_block2a2.port_a_logical_ram_depth = 64;
defparam ram_block2a2.port_a_logical_ram_width = 8;
defparam ram_block2a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_address_clear = "none";
defparam ram_block2a2.port_b_address_clock = "clock1";
defparam ram_block2a2.port_b_address_width = 6;
defparam ram_block2a2.port_b_data_out_clear = "none";
defparam ram_block2a2.port_b_data_out_clock = "none";
defparam ram_block2a2.port_b_data_width = 1;
defparam ram_block2a2.port_b_first_address = 0;
defparam ram_block2a2.port_b_first_bit_number = 2;
defparam ram_block2a2.port_b_last_address = 63;
defparam ram_block2a2.port_b_logical_ram_depth = 64;
defparam ram_block2a2.port_b_logical_ram_width = 8;
defparam ram_block2a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_read_enable_clock = "clock1";
defparam ram_block2a2.ram_block_type = "auto";

cycloneive_ram_block ram_block2a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a3_PORTBDATAOUT_bus));
defparam ram_block2a3.clk0_core_clock_enable = "ena0";
defparam ram_block2a3.clk1_core_clock_enable = "ena1";
defparam ram_block2a3.clk1_input_clock_enable = "ena1";
defparam ram_block2a3.data_interleave_offset_in_bits = 1;
defparam ram_block2a3.data_interleave_width_in_bits = 1;
defparam ram_block2a3.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a3.operation_mode = "dual_port";
defparam ram_block2a3.port_a_address_clear = "none";
defparam ram_block2a3.port_a_address_width = 6;
defparam ram_block2a3.port_a_data_out_clear = "none";
defparam ram_block2a3.port_a_data_out_clock = "none";
defparam ram_block2a3.port_a_data_width = 1;
defparam ram_block2a3.port_a_first_address = 0;
defparam ram_block2a3.port_a_first_bit_number = 3;
defparam ram_block2a3.port_a_last_address = 63;
defparam ram_block2a3.port_a_logical_ram_depth = 64;
defparam ram_block2a3.port_a_logical_ram_width = 8;
defparam ram_block2a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_address_clear = "none";
defparam ram_block2a3.port_b_address_clock = "clock1";
defparam ram_block2a3.port_b_address_width = 6;
defparam ram_block2a3.port_b_data_out_clear = "none";
defparam ram_block2a3.port_b_data_out_clock = "none";
defparam ram_block2a3.port_b_data_width = 1;
defparam ram_block2a3.port_b_first_address = 0;
defparam ram_block2a3.port_b_first_bit_number = 3;
defparam ram_block2a3.port_b_last_address = 63;
defparam ram_block2a3.port_b_logical_ram_depth = 64;
defparam ram_block2a3.port_b_logical_ram_width = 8;
defparam ram_block2a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_read_enable_clock = "clock1";
defparam ram_block2a3.ram_block_type = "auto";

cycloneive_ram_block ram_block2a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a4_PORTBDATAOUT_bus));
defparam ram_block2a4.clk0_core_clock_enable = "ena0";
defparam ram_block2a4.clk1_core_clock_enable = "ena1";
defparam ram_block2a4.clk1_input_clock_enable = "ena1";
defparam ram_block2a4.data_interleave_offset_in_bits = 1;
defparam ram_block2a4.data_interleave_width_in_bits = 1;
defparam ram_block2a4.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a4.operation_mode = "dual_port";
defparam ram_block2a4.port_a_address_clear = "none";
defparam ram_block2a4.port_a_address_width = 6;
defparam ram_block2a4.port_a_data_out_clear = "none";
defparam ram_block2a4.port_a_data_out_clock = "none";
defparam ram_block2a4.port_a_data_width = 1;
defparam ram_block2a4.port_a_first_address = 0;
defparam ram_block2a4.port_a_first_bit_number = 4;
defparam ram_block2a4.port_a_last_address = 63;
defparam ram_block2a4.port_a_logical_ram_depth = 64;
defparam ram_block2a4.port_a_logical_ram_width = 8;
defparam ram_block2a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_address_clear = "none";
defparam ram_block2a4.port_b_address_clock = "clock1";
defparam ram_block2a4.port_b_address_width = 6;
defparam ram_block2a4.port_b_data_out_clear = "none";
defparam ram_block2a4.port_b_data_out_clock = "none";
defparam ram_block2a4.port_b_data_width = 1;
defparam ram_block2a4.port_b_first_address = 0;
defparam ram_block2a4.port_b_first_bit_number = 4;
defparam ram_block2a4.port_b_last_address = 63;
defparam ram_block2a4.port_b_logical_ram_depth = 64;
defparam ram_block2a4.port_b_logical_ram_width = 8;
defparam ram_block2a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_read_enable_clock = "clock1";
defparam ram_block2a4.ram_block_type = "auto";

cycloneive_ram_block ram_block2a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a5_PORTBDATAOUT_bus));
defparam ram_block2a5.clk0_core_clock_enable = "ena0";
defparam ram_block2a5.clk1_core_clock_enable = "ena1";
defparam ram_block2a5.clk1_input_clock_enable = "ena1";
defparam ram_block2a5.data_interleave_offset_in_bits = 1;
defparam ram_block2a5.data_interleave_width_in_bits = 1;
defparam ram_block2a5.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a5.operation_mode = "dual_port";
defparam ram_block2a5.port_a_address_clear = "none";
defparam ram_block2a5.port_a_address_width = 6;
defparam ram_block2a5.port_a_data_out_clear = "none";
defparam ram_block2a5.port_a_data_out_clock = "none";
defparam ram_block2a5.port_a_data_width = 1;
defparam ram_block2a5.port_a_first_address = 0;
defparam ram_block2a5.port_a_first_bit_number = 5;
defparam ram_block2a5.port_a_last_address = 63;
defparam ram_block2a5.port_a_logical_ram_depth = 64;
defparam ram_block2a5.port_a_logical_ram_width = 8;
defparam ram_block2a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_address_clear = "none";
defparam ram_block2a5.port_b_address_clock = "clock1";
defparam ram_block2a5.port_b_address_width = 6;
defparam ram_block2a5.port_b_data_out_clear = "none";
defparam ram_block2a5.port_b_data_out_clock = "none";
defparam ram_block2a5.port_b_data_width = 1;
defparam ram_block2a5.port_b_first_address = 0;
defparam ram_block2a5.port_b_first_bit_number = 5;
defparam ram_block2a5.port_b_last_address = 63;
defparam ram_block2a5.port_b_logical_ram_depth = 64;
defparam ram_block2a5.port_b_logical_ram_width = 8;
defparam ram_block2a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_read_enable_clock = "clock1";
defparam ram_block2a5.ram_block_type = "auto";

cycloneive_ram_block ram_block2a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a6_PORTBDATAOUT_bus));
defparam ram_block2a6.clk0_core_clock_enable = "ena0";
defparam ram_block2a6.clk1_core_clock_enable = "ena1";
defparam ram_block2a6.clk1_input_clock_enable = "ena1";
defparam ram_block2a6.data_interleave_offset_in_bits = 1;
defparam ram_block2a6.data_interleave_width_in_bits = 1;
defparam ram_block2a6.logical_ram_name = "usb_system_jtag_uart:jtag_uart|usb_system_jtag_uart_scfifo_w:the_usb_system_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a6.operation_mode = "dual_port";
defparam ram_block2a6.port_a_address_clear = "none";
defparam ram_block2a6.port_a_address_width = 6;
defparam ram_block2a6.port_a_data_out_clear = "none";
defparam ram_block2a6.port_a_data_out_clock = "none";
defparam ram_block2a6.port_a_data_width = 1;
defparam ram_block2a6.port_a_first_address = 0;
defparam ram_block2a6.port_a_first_bit_number = 6;
defparam ram_block2a6.port_a_last_address = 63;
defparam ram_block2a6.port_a_logical_ram_depth = 64;
defparam ram_block2a6.port_a_logical_ram_width = 8;
defparam ram_block2a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_address_clear = "none";
defparam ram_block2a6.port_b_address_clock = "clock1";
defparam ram_block2a6.port_b_address_width = 6;
defparam ram_block2a6.port_b_data_out_clear = "none";
defparam ram_block2a6.port_b_data_out_clock = "none";
defparam ram_block2a6.port_b_data_width = 1;
defparam ram_block2a6.port_b_first_address = 0;
defparam ram_block2a6.port_b_first_bit_number = 6;
defparam ram_block2a6.port_b_last_address = 63;
defparam ram_block2a6.port_b_logical_ram_depth = 64;
defparam ram_block2a6.port_b_logical_ram_width = 8;
defparam ram_block2a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_read_enable_clock = "clock1";
defparam ram_block2a6.ram_block_type = "auto";

endmodule

module usb_system_usb_system_keycode (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	writedata,
	reset_n,
	Equal6,
	mem_used_1,
	always0,
	d_write,
	write_accepted,
	always01,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	[31:0] writedata;
input 	reset_n;
input 	Equal6;
input 	mem_used_1;
output 	always0;
input 	d_write;
input 	write_accepted;
output 	always01;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~2_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(Equal6),
	.datab(mem_used_1),
	.datac(W_alu_result_4),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hBFFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~1 (
	.dataa(d_write),
	.datab(W_alu_result_2),
	.datac(W_alu_result_3),
	.datad(write_accepted),
	.cin(gnd),
	.combout(always01),
	.cout());
defparam \always0~1 .lut_mask = 16'hBFFF;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAFFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAFFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAFFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAFFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAFFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAFFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAFFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAFFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~2 (
	.dataa(always0),
	.datab(always01),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hEFFF;
defparam \always0~2 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_keycode_1 (
	W_alu_result_7,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	writedata,
	Equal3,
	always0,
	reset_n,
	mem_used_1,
	always01,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	[31:0] writedata;
input 	Equal3;
input 	always0;
input 	reset_n;
input 	mem_used_1;
output 	always01;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~2_combout ;
wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cycloneive_lcell_comb \always0~1 (
	.dataa(W_alu_result_4),
	.datab(mem_used_1),
	.datac(Equal3),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(always01),
	.cout());
defparam \always0~1 .lut_mask = 16'hFFFB;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAFFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAFFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAFFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAFFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAFFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAFFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAFFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAFFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~2 (
	.dataa(always0),
	.datab(always01),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hEFFF;
defparam \always0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hBBBB;
defparam \always0~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0 (
	wire_pll7_clk_0,
	W_alu_result_7,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_8,
	W_alu_result_6,
	W_alu_result_24,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_5,
	readdata_6,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	Equal3,
	Equal6,
	mem_used_1,
	always0,
	d_write,
	write_accepted,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	altera_reset_synchronizer_int_chain_out,
	mem_used_11,
	always01,
	wait_latency_counter_11,
	wait_latency_counter_01,
	mem_used_12,
	always02,
	wait_latency_counter_12,
	wait_latency_counter_02,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	entries_1,
	entries_0,
	altera_reset_synchronizer_int_chain_out1,
	sink_in_reset,
	d_read,
	read_accepted,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	out_valid,
	src0_valid,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	mem_86_0,
	mem_68_0,
	src0_valid1,
	read_latency_shift_reg_04,
	read_latency_shift_reg_05,
	WideOr1,
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	src0_valid2,
	mem_67_04,
	mem_67_05,
	mem_67_06,
	mem_67_07,
	mem_67_08,
	out_valid1,
	out_data_buffer_67,
	av_ld_getting_data,
	waitrequest,
	mem_used_13,
	uav_write,
	mem_used_14,
	full,
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_5,
	F_pc_6,
	F_pc_4,
	F_pc_1,
	F_pc_3,
	i_read,
	F_pc_2,
	mem_used_15,
	av_waitrequest,
	Equal9,
	cpu_data_master_waitrequest,
	s0_cmd_valid,
	WideOr11,
	F_pc_0,
	src_data_38,
	mem,
	src_data_39,
	last_cycle,
	saved_grant_1,
	WideOr12,
	src_payload,
	src_data_68,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	src_data_61,
	src_data_60,
	src_data_381,
	src_data_391,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	out_data_buffer_32,
	out_data_buffer_321,
	out_data_buffer_33,
	out_data_buffer_331,
	out_data_buffer_34,
	out_data_buffer_341,
	out_data_buffer_35,
	out_data_buffer_351,
	sink_ready,
	WideOr13,
	local_read,
	mem1,
	m0_write,
	src1_valid,
	src_payload1,
	out_valid2,
	src_payload2,
	WideOr14,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	hbreak_enabled,
	out_data_buffer_0,
	av_readdata_pre_0,
	av_readdata_pre_01,
	out_data_buffer_1,
	av_readdata_pre_1,
	av_readdata_pre_11,
	out_data_buffer_2,
	av_readdata_pre_2,
	av_readdata_pre_30,
	src_payload3,
	av_readdata_pre_3,
	out_data_buffer_4,
	av_readdata_pre_4,
	out_payload_0,
	src_data_0,
	out_data_buffer_22,
	av_readdata_pre_22,
	av_readdata_pre_23,
	out_data_buffer_23,
	out_data_buffer_24,
	av_readdata_pre_24,
	av_readdata_pre_25,
	out_data_buffer_25,
	out_data_buffer_26,
	av_readdata_pre_26,
	out_data_buffer_11,
	av_readdata_pre_111,
	out_data_buffer_13,
	av_readdata_pre_13,
	src_payload4,
	av_readdata_pre_16,
	av_readdata_pre_12,
	out_data_buffer_12,
	out_data_buffer_5,
	av_readdata_pre_5,
	out_data_buffer_14,
	av_readdata_pre_14,
	out_data_buffer_15,
	av_readdata_pre_15,
	av_readdata_pre_10,
	out_data_buffer_10,
	out_data_buffer_9,
	av_readdata_pre_9,
	out_data_buffer_8,
	av_readdata_pre_8,
	out_data_buffer_7,
	av_readdata_pre_7,
	out_data_buffer_6,
	av_readdata_pre_6,
	src_payload5,
	av_readdata_pre_20,
	out_data_buffer_18,
	av_readdata_pre_18,
	out_data_buffer_19,
	av_readdata_pre_19,
	out_data_buffer_17,
	av_readdata_pre_17,
	src_payload6,
	av_readdata_pre_21,
	av_readdata_pre_27,
	out_data_buffer_27,
	out_data_buffer_28,
	av_readdata_pre_28,
	av_readdata_pre_31,
	out_data_buffer_31,
	out_data_buffer_30,
	av_readdata_pre_301,
	av_readdata_pre_29,
	out_data_buffer_29,
	mem2,
	src_data_461,
	out_payload_1,
	src_data_1,
	src_payload7,
	out_payload_2,
	src_data_2,
	src_data_3,
	out_payload_3,
	src_data_31,
	out_payload_4,
	src_data_4,
	out_payload_5,
	src_data_5,
	out_payload_6,
	src_data_6,
	out_payload_7,
	src_data_7,
	out_payload_8,
	src_data_8,
	av_readdata_9,
	av_readdata_8,
	readdata_01,
	readdata_11,
	readdata_4,
	out_payload_9,
	src_data_9,
	out_payload_10,
	src_data_10,
	out_payload_11,
	src_data_11,
	out_payload_12,
	src_data_12,
	out_payload_13,
	src_data_13,
	out_payload_14,
	src_data_14,
	out_payload_15,
	src_data_15,
	src_data_16,
	src_data_17,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	b_full,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	read_0,
	av_readdata_0,
	readdata_02,
	readdata_03,
	readdata_04,
	readdata_05,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_111,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_14,
	readdata_15,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_20,
	readdata_18,
	readdata_19,
	readdata_17,
	src_payload40,
	readdata_21,
	src_payload41,
	readdata_27,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	out_data_buffer_241,
	readdata_28,
	out_data_buffer_281,
	out_data_buffer_271,
	readdata_31,
	out_data_buffer_261,
	readdata_30,
	out_data_buffer_251,
	readdata_29,
	av_readdata_1,
	readdata_110,
	readdata_112,
	readdata_113,
	readdata_114,
	av_readdata_2,
	readdata_210,
	readdata_211,
	readdata_212,
	readdata_213,
	readdata_32,
	readdata_33,
	av_readdata_3,
	readdata_34,
	readdata_35,
	av_readdata_4,
	readdata_41,
	readdata_42,
	readdata_43,
	readdata_44,
	av_readdata_5,
	readdata_51,
	readdata_52,
	readdata_53,
	readdata_54,
	av_readdata_6,
	readdata_61,
	readdata_62,
	readdata_63,
	readdata_64,
	av_readdata_7,
	readdata_71,
	readdata_72,
	readdata_73,
	readdata_74,
	readdata_81,
	readdata_82,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_01,
	counter_reg_bit_11,
	counter_reg_bit_41,
	counter_reg_bit_51,
	readdata_91,
	readdata_92,
	ac,
	readdata_101,
	readdata_102,
	readdata_115,
	readdata_116,
	readdata_121,
	readdata_122,
	readdata_131,
	readdata_132,
	woverflow,
	readdata_141,
	readdata_142,
	readdata_151,
	readdata_152,
	rvalid,
	readdata_161,
	readdata_162,
	readdata_171,
	readdata_172,
	src_payload46,
	src_payload47,
	src_data_382,
	src_data_392,
	src_data_401,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_32,
	out_data_buffer_311,
	out_data_buffer_301,
	out_data_buffer_291,
	src_payload48,
	src_payload49,
	src_payload50,
	za_valid,
	src_payload51,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	src_payload52,
	src_payload53,
	src_payload54,
	src_data_34,
	src_payload55,
	src_payload56,
	src_payload57,
	src_data_35,
	src_payload58,
	src_payload59,
	src_payload60,
	src_data_33,
	src_payload61,
	src_payload62,
	src_payload63,
	src_payload64,
	src_payload65,
	src_payload66,
	src_payload67,
	src_payload68,
	src_payload69,
	src_payload70,
	src_payload71,
	src_payload72,
	src_payload73,
	src_payload74,
	src_payload75,
	src_payload76,
	src_payload77,
	src_payload78,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_22,
	za_data_23,
	za_data_24,
	za_data_25,
	za_data_26,
	za_data_11,
	za_data_13,
	za_data_16,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_10,
	za_data_9,
	za_data_8,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_18,
	za_data_19,
	za_data_17,
	za_data_21,
	za_data_27,
	za_data_28,
	za_data_31,
	za_data_30,
	za_data_29,
	m0_write1,
	m0_read,
	m0_write2,
	src_data_21,
	src_data_410,
	src_data_510,
	src_data_63,
	src_data_71,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_7;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_8;
input 	W_alu_result_6;
input 	W_alu_result_24;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_28;
input 	W_alu_result_27;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	readdata_0;
input 	readdata_1;
input 	readdata_2;
input 	readdata_3;
input 	readdata_5;
input 	readdata_6;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
output 	Equal3;
output 	Equal6;
output 	mem_used_1;
input 	always0;
input 	d_write;
output 	write_accepted;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	altera_reset_synchronizer_int_chain_out;
output 	mem_used_11;
input 	always01;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
output 	mem_used_12;
input 	always02;
output 	wait_latency_counter_12;
output 	wait_latency_counter_02;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	entries_1;
input 	entries_0;
input 	altera_reset_synchronizer_int_chain_out1;
input 	sink_in_reset;
input 	d_read;
output 	read_accepted;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg_01;
input 	out_valid;
output 	src0_valid;
output 	read_latency_shift_reg_02;
output 	read_latency_shift_reg_03;
output 	mem_86_0;
output 	mem_68_0;
output 	src0_valid1;
output 	read_latency_shift_reg_04;
output 	read_latency_shift_reg_05;
output 	WideOr1;
output 	mem_67_0;
output 	mem_67_01;
output 	mem_67_02;
output 	mem_67_03;
output 	src0_valid2;
output 	mem_67_04;
output 	mem_67_05;
output 	mem_67_06;
output 	mem_67_07;
output 	mem_67_08;
output 	out_valid1;
output 	out_data_buffer_67;
input 	av_ld_getting_data;
input 	waitrequest;
output 	mem_used_13;
output 	uav_write;
output 	mem_used_14;
input 	full;
input 	F_pc_26;
input 	F_pc_25;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_4;
input 	F_pc_1;
input 	F_pc_3;
input 	i_read;
input 	F_pc_2;
output 	mem_used_15;
input 	av_waitrequest;
output 	Equal9;
output 	cpu_data_master_waitrequest;
input 	s0_cmd_valid;
output 	WideOr11;
input 	F_pc_0;
output 	src_data_38;
output 	mem;
output 	src_data_39;
output 	last_cycle;
output 	saved_grant_1;
output 	WideOr12;
output 	src_payload;
output 	src_data_68;
output 	src_data_48;
output 	src_data_62;
output 	src_data_49;
output 	src_data_51;
output 	src_data_50;
output 	src_data_53;
output 	src_data_52;
output 	src_data_55;
output 	src_data_54;
output 	src_data_57;
output 	src_data_56;
output 	src_data_59;
output 	src_data_58;
output 	src_data_61;
output 	src_data_60;
output 	src_data_381;
output 	src_data_391;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	out_data_buffer_32;
output 	out_data_buffer_321;
output 	out_data_buffer_33;
output 	out_data_buffer_331;
output 	out_data_buffer_34;
output 	out_data_buffer_341;
output 	out_data_buffer_35;
output 	out_data_buffer_351;
output 	sink_ready;
output 	WideOr13;
output 	local_read;
output 	mem1;
output 	m0_write;
output 	src1_valid;
output 	src_payload1;
output 	out_valid2;
output 	src_payload2;
output 	WideOr14;
output 	av_readdatavalid;
output 	av_readdatavalid1;
output 	av_readdatavalid2;
input 	hbreak_enabled;
output 	out_data_buffer_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_01;
output 	out_data_buffer_1;
output 	av_readdata_pre_1;
output 	av_readdata_pre_11;
output 	out_data_buffer_2;
output 	av_readdata_pre_2;
output 	av_readdata_pre_30;
output 	src_payload3;
output 	av_readdata_pre_3;
output 	out_data_buffer_4;
output 	av_readdata_pre_4;
input 	out_payload_0;
output 	src_data_0;
output 	out_data_buffer_22;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	av_readdata_pre_26;
output 	out_data_buffer_11;
output 	av_readdata_pre_111;
output 	out_data_buffer_13;
output 	av_readdata_pre_13;
output 	src_payload4;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	av_readdata_pre_5;
output 	out_data_buffer_14;
output 	av_readdata_pre_14;
output 	out_data_buffer_15;
output 	av_readdata_pre_15;
output 	av_readdata_pre_10;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	av_readdata_pre_9;
output 	out_data_buffer_8;
output 	av_readdata_pre_8;
output 	out_data_buffer_7;
output 	av_readdata_pre_7;
output 	out_data_buffer_6;
output 	av_readdata_pre_6;
output 	src_payload5;
output 	av_readdata_pre_20;
output 	out_data_buffer_18;
output 	av_readdata_pre_18;
output 	out_data_buffer_19;
output 	av_readdata_pre_19;
output 	out_data_buffer_17;
output 	av_readdata_pre_17;
output 	src_payload6;
output 	av_readdata_pre_21;
output 	av_readdata_pre_27;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	av_readdata_pre_28;
output 	av_readdata_pre_31;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	av_readdata_pre_301;
output 	av_readdata_pre_29;
output 	out_data_buffer_29;
output 	mem2;
output 	src_data_461;
input 	out_payload_1;
output 	src_data_1;
output 	src_payload7;
input 	out_payload_2;
output 	src_data_2;
output 	src_data_3;
input 	out_payload_3;
output 	src_data_31;
input 	out_payload_4;
output 	src_data_4;
input 	out_payload_5;
output 	src_data_5;
input 	out_payload_6;
output 	src_data_6;
input 	out_payload_7;
output 	src_data_7;
input 	out_payload_8;
output 	src_data_8;
input 	av_readdata_9;
input 	av_readdata_8;
input 	readdata_01;
input 	readdata_11;
input 	readdata_4;
input 	out_payload_9;
output 	src_data_9;
input 	out_payload_10;
output 	src_data_10;
input 	out_payload_11;
output 	src_data_11;
input 	out_payload_12;
output 	src_data_12;
input 	out_payload_13;
output 	src_data_13;
input 	out_payload_14;
output 	src_data_14;
input 	out_payload_15;
output 	src_data_15;
output 	src_data_16;
output 	src_data_17;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
input 	b_full;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
output 	src_payload35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
input 	read_0;
input 	av_readdata_0;
input 	readdata_02;
input 	readdata_03;
input 	readdata_04;
input 	readdata_05;
input 	readdata_22;
input 	readdata_23;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_111;
input 	readdata_13;
input 	readdata_16;
input 	readdata_12;
input 	readdata_14;
input 	readdata_15;
input 	readdata_10;
input 	readdata_9;
input 	readdata_8;
input 	readdata_7;
input 	readdata_20;
input 	readdata_18;
input 	readdata_19;
input 	readdata_17;
output 	src_payload40;
input 	readdata_21;
output 	src_payload41;
input 	readdata_27;
output 	src_payload42;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	out_data_buffer_241;
input 	readdata_28;
output 	out_data_buffer_281;
output 	out_data_buffer_271;
input 	readdata_31;
output 	out_data_buffer_261;
input 	readdata_30;
output 	out_data_buffer_251;
input 	readdata_29;
input 	av_readdata_1;
input 	readdata_110;
input 	readdata_112;
input 	readdata_113;
input 	readdata_114;
input 	av_readdata_2;
input 	readdata_210;
input 	readdata_211;
input 	readdata_212;
input 	readdata_213;
input 	readdata_32;
input 	readdata_33;
input 	av_readdata_3;
input 	readdata_34;
input 	readdata_35;
input 	av_readdata_4;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
input 	readdata_44;
input 	av_readdata_5;
input 	readdata_51;
input 	readdata_52;
input 	readdata_53;
input 	readdata_54;
input 	av_readdata_6;
input 	readdata_61;
input 	readdata_62;
input 	readdata_63;
input 	readdata_64;
input 	av_readdata_7;
input 	readdata_71;
input 	readdata_72;
input 	readdata_73;
input 	readdata_74;
input 	readdata_81;
input 	readdata_82;
input 	counter_reg_bit_3;
input 	counter_reg_bit_0;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	b_full1;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	b_non_empty;
input 	counter_reg_bit_31;
input 	counter_reg_bit_21;
input 	counter_reg_bit_01;
input 	counter_reg_bit_11;
input 	counter_reg_bit_41;
input 	counter_reg_bit_51;
input 	readdata_91;
input 	readdata_92;
input 	ac;
input 	readdata_101;
input 	readdata_102;
input 	readdata_115;
input 	readdata_116;
input 	readdata_121;
input 	readdata_122;
input 	readdata_131;
input 	readdata_132;
input 	woverflow;
input 	readdata_141;
input 	readdata_142;
input 	readdata_151;
input 	readdata_152;
input 	rvalid;
input 	readdata_161;
input 	readdata_162;
input 	readdata_171;
input 	readdata_172;
output 	src_payload46;
output 	src_payload47;
output 	src_data_382;
output 	src_data_392;
output 	src_data_401;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_32;
output 	out_data_buffer_311;
output 	out_data_buffer_301;
output 	out_data_buffer_291;
output 	src_payload48;
output 	src_payload49;
output 	src_payload50;
input 	za_valid;
output 	src_payload51;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
output 	src_payload52;
output 	src_payload53;
output 	src_payload54;
output 	src_data_34;
output 	src_payload55;
output 	src_payload56;
output 	src_payload57;
output 	src_data_35;
output 	src_payload58;
output 	src_payload59;
output 	src_payload60;
output 	src_data_33;
output 	src_payload61;
output 	src_payload62;
output 	src_payload63;
output 	src_payload64;
output 	src_payload65;
output 	src_payload66;
output 	src_payload67;
output 	src_payload68;
output 	src_payload69;
output 	src_payload70;
output 	src_payload71;
output 	src_payload72;
output 	src_payload73;
output 	src_payload74;
output 	src_payload75;
output 	src_payload76;
output 	src_payload77;
output 	src_payload78;
input 	za_data_0;
input 	za_data_1;
input 	za_data_2;
input 	za_data_3;
input 	za_data_4;
input 	za_data_22;
input 	za_data_23;
input 	za_data_24;
input 	za_data_25;
input 	za_data_26;
input 	za_data_11;
input 	za_data_13;
input 	za_data_16;
input 	za_data_12;
input 	za_data_5;
input 	za_data_14;
input 	za_data_15;
input 	za_data_10;
input 	za_data_9;
input 	za_data_8;
input 	za_data_7;
input 	za_data_6;
input 	za_data_20;
input 	za_data_18;
input 	za_data_19;
input 	za_data_17;
input 	za_data_21;
input 	za_data_27;
input 	za_data_28;
input 	za_data_31;
input 	za_data_30;
input 	za_data_29;
output 	m0_write1;
output 	m0_read;
output 	m0_write2;
output 	src_data_21;
output 	src_data_410;
output 	src_data_510;
output 	src_data_63;
output 	src_data_71;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \router|Equal1~0_combout ;
wire \keycode_s1_translator|read_latency_shift_reg~2_combout ;
wire \keycode_s1_translator|read_latency_shift_reg~3_combout ;
wire \sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \clocks_pll_slave_translator|read_latency_shift_reg[0]~q ;
wire \clocks_pll_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \clocks_pll_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \crosser_002|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_002|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \router|Equal2~5_combout ;
wire \cmd_mux_002|saved_grant[0]~q ;
wire \router|always1~2_combout ;
wire \all_switches_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \all_switches_s1_translator|wait_latency_counter[1]~1_combout ;
wire \all_switches_s1_translator|waitrequest_reset_override~q ;
wire \cmd_mux_003|saved_grant[0]~q ;
wire \clock_crossing_io_s0_agent_rsp_fifo|mem_used[128]~q ;
wire \router|Equal1~2_combout ;
wire \cmd_mux_001|saved_grant[0]~q ;
wire \cpu_data_master_translator|uav_read~0_combout ;
wire \router|always1~3_combout ;
wire \cmd_demux|sink_ready~2_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \router_001|Equal1~4_combout ;
wire \router_001|Equal2~1_combout ;
wire \cpu_instruction_master_translator|read_accepted~q ;
wire \router_001|always1~1_combout ;
wire \cmd_mux_001|src_valid~0_combout ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \sysid_qsys_0_control_slave_agent|m0_write~0_combout ;
wire \sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ;
wire \sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ;
wire \router|Equal9~0_combout ;
wire \cmd_demux|sink_ready~7_combout ;
wire \crosser|clock_xer|in_data_toggle~q ;
wire \crosser|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \router|always1~4_combout ;
wire \red_leds_s1_translator|wait_latency_counter[1]~1_combout ;
wire \led_s1_translator|wait_latency_counter[0]~1_combout ;
wire \cmd_demux|WideOr0~7_combout ;
wire \router|Equal5~0_combout ;
wire \router|Equal3~6_combout ;
wire \cpu_instruction_master_translator|uav_read~0_combout ;
wire \cmd_mux_003|saved_grant[1]~q ;
wire \router_001|Equal2~2_combout ;
wire \router|Equal7~0_combout ;
wire \sdram_s1_agent_rsp_fifo|mem_used[7]~q ;
wire \cmd_mux_006|saved_grant[0]~q ;
wire \crosser_001|clock_xer|out_valid~combout ;
wire \crosser|clock_xer|out_data_toggle_flopped~q ;
wire \crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser|clock_xer|out_valid~combout ;
wire \crosser|clock_xer|out_data_buffer[67]~q ;
wire \crosser_001|clock_xer|out_data_buffer[68]~q ;
wire \crosser|clock_xer|out_data_buffer[68]~q ;
wire \crosser_001|clock_xer|out_data_buffer[48]~q ;
wire \crosser|clock_xer|out_data_buffer[48]~q ;
wire \crosser_001|clock_xer|out_data_buffer[62]~q ;
wire \crosser|clock_xer|out_data_buffer[62]~q ;
wire \crosser_001|clock_xer|out_data_buffer[49]~q ;
wire \crosser|clock_xer|out_data_buffer[49]~q ;
wire \crosser_001|clock_xer|out_data_buffer[51]~q ;
wire \crosser|clock_xer|out_data_buffer[51]~q ;
wire \crosser_001|clock_xer|out_data_buffer[50]~q ;
wire \crosser|clock_xer|out_data_buffer[50]~q ;
wire \crosser_001|clock_xer|out_data_buffer[53]~q ;
wire \crosser|clock_xer|out_data_buffer[53]~q ;
wire \crosser_001|clock_xer|out_data_buffer[52]~q ;
wire \crosser|clock_xer|out_data_buffer[52]~q ;
wire \crosser_001|clock_xer|out_data_buffer[55]~q ;
wire \crosser|clock_xer|out_data_buffer[55]~q ;
wire \crosser_001|clock_xer|out_data_buffer[54]~q ;
wire \crosser|clock_xer|out_data_buffer[54]~q ;
wire \crosser_001|clock_xer|out_data_buffer[57]~q ;
wire \crosser|clock_xer|out_data_buffer[57]~q ;
wire \crosser_001|clock_xer|out_data_buffer[56]~q ;
wire \crosser|clock_xer|out_data_buffer[56]~q ;
wire \crosser_001|clock_xer|out_data_buffer[59]~q ;
wire \crosser|clock_xer|out_data_buffer[59]~q ;
wire \crosser_001|clock_xer|out_data_buffer[58]~q ;
wire \crosser|clock_xer|out_data_buffer[58]~q ;
wire \crosser_001|clock_xer|out_data_buffer[61]~q ;
wire \crosser|clock_xer|out_data_buffer[61]~q ;
wire \crosser_001|clock_xer|out_data_buffer[60]~q ;
wire \crosser|clock_xer|out_data_buffer[60]~q ;
wire \crosser_001|clock_xer|out_data_buffer[38]~q ;
wire \crosser|clock_xer|out_data_buffer[38]~q ;
wire \crosser_001|clock_xer|out_data_buffer[39]~q ;
wire \crosser|clock_xer|out_data_buffer[39]~q ;
wire \crosser_001|clock_xer|out_data_buffer[40]~q ;
wire \crosser|clock_xer|out_data_buffer[40]~q ;
wire \crosser_001|clock_xer|out_data_buffer[41]~q ;
wire \crosser|clock_xer|out_data_buffer[41]~q ;
wire \crosser_001|clock_xer|out_data_buffer[42]~q ;
wire \crosser|clock_xer|out_data_buffer[42]~q ;
wire \crosser_001|clock_xer|out_data_buffer[43]~q ;
wire \crosser|clock_xer|out_data_buffer[43]~q ;
wire \crosser_001|clock_xer|out_data_buffer[44]~q ;
wire \crosser|clock_xer|out_data_buffer[44]~q ;
wire \crosser_001|clock_xer|out_data_buffer[45]~q ;
wire \crosser|clock_xer|out_data_buffer[45]~q ;
wire \crosser_001|clock_xer|out_data_buffer[46]~q ;
wire \crosser|clock_xer|out_data_buffer[46]~q ;
wire \crosser_001|clock_xer|out_data_buffer[47]~q ;
wire \crosser|clock_xer|out_data_buffer[47]~q ;
wire \router|Equal6~2_combout ;
wire \red_leds_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_mux_001|src_data[68]~combout ;
wire \router_001|always1~2_combout ;
wire \sysid_qsys_0_control_slave_translator|read_latency_shift_reg~1_combout ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \cpu_debug_mem_slave_agent_rsp_fifo|mem~0_combout ;
wire \clocks_pll_slave_translator|read_latency_shift_reg~0_combout ;
wire \led_s1_translator|read_latency_shift_reg~0_combout ;
wire \router|always1~5_combout ;
wire \cmd_demux|sink_ready~12_combout ;
wire \all_switches_s1_agent|m0_write~0_combout ;
wire \cmd_demux|sink_ready~13_combout ;
wire \cmd_demux_001|src2_valid~0_combout ;
wire \router|Equal1~3_combout ;
wire \router|always1~6_combout ;
wire \cmd_mux_001|WideOr1~combout ;
wire \sysid_qsys_0_control_slave_agent|cp_ready~0_combout ;
wire \crosser_003|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_003|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser_003|clock_xer|out_data_buffer[67]~q ;
wire \router_001|Equal1~5_combout ;
wire \crosser_001|clock_xer|take_in_data~2_combout ;
wire \cmd_mux_001|src_payload~0_combout ;
wire \cmd_demux|sink_ready~14_combout ;
wire \crosser_003|clock_xer|out_data_buffer[3]~q ;
wire \crosser_001|clock_xer|out_data_buffer[107]~q ;
wire \crosser|clock_xer|out_data_buffer[107]~q ;
wire \cmd_mux_006|src_payload[0]~combout ;
wire \crosser|clock_xer|out_data_buffer[66]~q ;
wire \sdram_s1_agent|nonposted_write_endofpacket~0_combout ;
wire \sdram_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \sdram_s1_agent_rdata_fifo|out_valid~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][86]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \crosser_003|clock_xer|in_data_toggle~q ;
wire \crosser_003|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_002|clock_xer|in_data_toggle~q ;
wire \crosser_002|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \router_008|always0~0_combout ;
wire \rsp_demux_006|WideOr0~1_combout ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \led_s1_translator|av_readdata_pre[0]~q ;
wire \keycode_s1_translator|av_readdata_pre[0]~q ;
wire \all_switches_s1_translator|av_readdata_pre[0]~q ;
wire \red_leds_s1_translator|av_readdata_pre[0]~q ;
wire \crosser_002|clock_xer|out_data_buffer[0]~q ;
wire \crosser_003|clock_xer|out_data_buffer[16]~q ;
wire \crosser_003|clock_xer|out_data_buffer[20]~q ;
wire \crosser_003|clock_xer|out_data_buffer[21]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \crosser_002|clock_xer|take_in_data~0_combout ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \led_s1_translator|av_readdata_pre[1]~q ;
wire \keycode_s1_translator|av_readdata_pre[1]~q ;
wire \all_switches_s1_translator|av_readdata_pre[1]~q ;
wire \red_leds_s1_translator|av_readdata_pre[1]~q ;
wire \crosser_002|clock_xer|out_data_buffer[1]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \led_s1_translator|av_readdata_pre[2]~q ;
wire \keycode_s1_translator|av_readdata_pre[2]~q ;
wire \all_switches_s1_translator|av_readdata_pre[2]~q ;
wire \red_leds_s1_translator|av_readdata_pre[2]~q ;
wire \crosser_002|clock_xer|out_data_buffer[2]~q ;
wire \all_switches_s1_translator|av_readdata_pre[3]~q ;
wire \red_leds_s1_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \led_s1_translator|av_readdata_pre[3]~q ;
wire \keycode_s1_translator|av_readdata_pre[3]~q ;
wire \crosser_002|clock_xer|out_data_buffer[3]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \led_s1_translator|av_readdata_pre[4]~q ;
wire \keycode_s1_translator|av_readdata_pre[4]~q ;
wire \all_switches_s1_translator|av_readdata_pre[4]~q ;
wire \red_leds_s1_translator|av_readdata_pre[4]~q ;
wire \crosser_002|clock_xer|out_data_buffer[4]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \led_s1_translator|av_readdata_pre[5]~q ;
wire \keycode_s1_translator|av_readdata_pre[5]~q ;
wire \all_switches_s1_translator|av_readdata_pre[5]~q ;
wire \red_leds_s1_translator|av_readdata_pre[5]~q ;
wire \crosser_002|clock_xer|out_data_buffer[5]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \led_s1_translator|av_readdata_pre[6]~q ;
wire \keycode_s1_translator|av_readdata_pre[6]~q ;
wire \all_switches_s1_translator|av_readdata_pre[6]~q ;
wire \red_leds_s1_translator|av_readdata_pre[6]~q ;
wire \crosser_002|clock_xer|out_data_buffer[6]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \led_s1_translator|av_readdata_pre[7]~q ;
wire \keycode_s1_translator|av_readdata_pre[7]~q ;
wire \all_switches_s1_translator|av_readdata_pre[7]~q ;
wire \red_leds_s1_translator|av_readdata_pre[7]~q ;
wire \crosser_002|clock_xer|out_data_buffer[7]~q ;
wire \all_switches_s1_translator|av_readdata_pre[8]~q ;
wire \red_leds_s1_translator|av_readdata_pre[8]~q ;
wire \crosser_002|clock_xer|out_data_buffer[8]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \cmd_mux_001|src_data[38]~combout ;
wire \all_switches_s1_translator|av_readdata_pre[9]~q ;
wire \red_leds_s1_translator|av_readdata_pre[9]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \crosser_002|clock_xer|out_data_buffer[9]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \all_switches_s1_translator|av_readdata_pre[10]~q ;
wire \red_leds_s1_translator|av_readdata_pre[10]~q ;
wire \crosser_002|clock_xer|out_data_buffer[10]~q ;
wire \all_switches_s1_translator|av_readdata_pre[11]~q ;
wire \crosser_002|clock_xer|out_data_buffer[11]~q ;
wire \red_leds_s1_translator|av_readdata_pre[11]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \all_switches_s1_translator|av_readdata_pre[12]~q ;
wire \red_leds_s1_translator|av_readdata_pre[12]~q ;
wire \crosser_002|clock_xer|out_data_buffer[12]~q ;
wire \all_switches_s1_translator|av_readdata_pre[13]~q ;
wire \red_leds_s1_translator|av_readdata_pre[13]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \crosser_002|clock_xer|out_data_buffer[13]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \all_switches_s1_translator|av_readdata_pre[14]~q ;
wire \red_leds_s1_translator|av_readdata_pre[14]~q ;
wire \crosser_002|clock_xer|out_data_buffer[14]~q ;
wire \all_switches_s1_translator|av_readdata_pre[15]~q ;
wire \red_leds_s1_translator|av_readdata_pre[15]~q ;
wire \crosser_002|clock_xer|out_data_buffer[15]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \all_switches_s1_translator|av_readdata_pre[16]~q ;
wire \crosser_002|clock_xer|out_data_buffer[16]~q ;
wire \red_leds_s1_translator|av_readdata_pre[16]~q ;
wire \all_switches_s1_translator|av_readdata_pre[17]~q ;
wire \crosser_002|clock_xer|out_data_buffer[17]~q ;
wire \red_leds_s1_translator|av_readdata_pre[17]~q ;
wire \crosser_001|clock_xer|out_data_buffer[86]~q ;
wire \crosser|clock_xer|out_data_buffer[0]~q ;
wire \crosser|clock_xer|out_data_buffer[1]~q ;
wire \crosser|clock_xer|out_data_buffer[2]~q ;
wire \crosser|clock_xer|out_data_buffer[3]~q ;
wire \crosser|clock_xer|out_data_buffer[4]~q ;
wire \crosser|clock_xer|out_data_buffer[5]~q ;
wire \crosser|clock_xer|out_data_buffer[6]~q ;
wire \crosser|clock_xer|out_data_buffer[7]~q ;
wire \crosser|clock_xer|out_data_buffer[8]~q ;
wire \crosser|clock_xer|out_data_buffer[9]~q ;
wire \crosser|clock_xer|out_data_buffer[10]~q ;
wire \crosser|clock_xer|out_data_buffer[11]~q ;
wire \crosser|clock_xer|out_data_buffer[12]~q ;
wire \crosser|clock_xer|out_data_buffer[13]~q ;
wire \crosser|clock_xer|out_data_buffer[14]~q ;
wire \crosser|clock_xer|out_data_buffer[15]~q ;
wire \crosser|clock_xer|out_data_buffer[16]~q ;
wire \crosser|clock_xer|out_data_buffer[17]~q ;
wire \crosser|clock_xer|out_data_buffer[18]~q ;
wire \crosser|clock_xer|out_data_buffer[19]~q ;
wire \crosser|clock_xer|out_data_buffer[20]~q ;
wire \crosser|clock_xer|out_data_buffer[21]~q ;
wire \crosser|clock_xer|out_data_buffer[22]~q ;
wire \crosser|clock_xer|out_data_buffer[23]~q ;
wire \crosser|clock_xer|out_data_buffer[24]~q ;
wire \crosser|clock_xer|out_data_buffer[25]~q ;
wire \crosser|clock_xer|out_data_buffer[26]~q ;
wire \crosser|clock_xer|out_data_buffer[27]~q ;
wire \crosser|clock_xer|out_data_buffer[28]~q ;
wire \crosser|clock_xer|out_data_buffer[29]~q ;
wire \crosser|clock_xer|out_data_buffer[30]~q ;
wire \crosser|clock_xer|out_data_buffer[31]~q ;
wire \crosser_002|clock_xer|out_data_buffer[18]~q ;
wire \crosser_002|clock_xer|out_data_buffer[23]~q ;
wire \crosser_002|clock_xer|out_data_buffer[22]~q ;
wire \crosser_002|clock_xer|out_data_buffer[21]~q ;
wire \crosser_002|clock_xer|out_data_buffer[20]~q ;
wire \crosser_002|clock_xer|out_data_buffer[19]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[0]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[1]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[2]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[3]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[4]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[22]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[23]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[24]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[25]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[26]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[11]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[13]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[16]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[12]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[5]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[14]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[15]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[10]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[9]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[8]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[7]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[6]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[20]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[18]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[19]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[17]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[21]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[27]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[28]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[31]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[30]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[29]~q ;


usb_system_altera_avalon_sc_fifo_5 keycode_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_used_1(mem_used_1),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.read_latency_shift_reg(\keycode_s1_translator|read_latency_shift_reg~2_combout ),
	.read_latency_shift_reg1(\keycode_s1_translator|read_latency_shift_reg~3_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_67_0(mem_67_05),
	.clk(clk_clk));

usb_system_altera_avalon_sc_fifo_1 clock_crossing_io_s0_agent_rsp_fifo(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.sink_in_reset(sink_in_reset),
	.read_latency_shift_reg(\keycode_s1_translator|read_latency_shift_reg~3_combout ),
	.out_valid(out_valid),
	.mem_67_0(mem_67_02),
	.full(full),
	.mem_used_128(\clock_crossing_io_s0_agent_rsp_fifo|mem_used[128]~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.m0_write(m0_write),
	.clk(clk_clk));

usb_system_altera_merlin_slave_agent_1 clock_crossing_io_s0_agent(
	.W_alu_result_24(W_alu_result_24),
	.Equal1(\router|Equal1~0_combout ),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.mem_used_128(\clock_crossing_io_s0_agent_rsp_fifo|mem_used[128]~q ),
	.Equal11(\router|Equal1~3_combout ),
	.m0_write(m0_write),
	.m0_read(m0_read),
	.m0_write1(m0_write2));

usb_system_altera_avalon_sc_fifo_2 clocks_pll_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.sink_in_reset(sink_in_reset),
	.read_latency_shift_reg_0(\clocks_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\clocks_pll_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\clocks_pll_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(mem_67_04),
	.uav_write(uav_write),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(mem_used_14),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.uav_read1(\cpu_instruction_master_translator|uav_read~0_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.WideOr1(WideOr11),
	.mem(mem),
	.mem1(mem1),
	.read_latency_shift_reg(\clocks_pll_slave_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

usb_system_altera_avalon_sc_fifo_3 cpu_debug_mem_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_01),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_13),
	.uav_write(uav_write),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.uav_read1(\cpu_instruction_master_translator|uav_read~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.mem(\cpu_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.local_read(local_read),
	.mem1(mem2),
	.clk(clk_clk));

usb_system_altera_merlin_slave_agent_3 cpu_debug_mem_slave_agent(
	.WideOr1(WideOr13),
	.mem(\cpu_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.local_read(local_read));

usb_system_altera_avalon_sc_fifo_10 sysid_qsys_0_control_slave_agent_rsp_fifo(
	.reset(altera_reset_synchronizer_int_chain_out),
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(mem_67_0),
	.uav_write(uav_write),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.src_data_68(\cmd_mux_001|src_data[68]~combout ),
	.read_latency_shift_reg(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg~1_combout ),
	.WideOr1(\cmd_mux_001|WideOr1~combout ),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ),
	.clk(clk_clk));

usb_system_altera_merlin_slave_agent_9 sysid_qsys_0_control_slave_agent(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\sysid_qsys_0_control_slave_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ));

usb_system_altera_avalon_sc_fifo_4 jtag_uart_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.mem_67_0(mem_67_03),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.mem_used_1(mem_used_15),
	.av_waitrequest(av_waitrequest),
	.Equal9(Equal9),
	.sink_ready(sink_ready),
	.clk(clk_clk));

usb_system_altera_merlin_master_agent_1 cpu_instruction_master_agent(
	.mem_67_0(mem_67_0),
	.mem_67_01(mem_67_01),
	.mem_67_02(mem_67_04),
	.src1_valid(src1_valid),
	.src_payload(src_payload1),
	.out_valid(out_valid2),
	.src_payload1(src_payload2),
	.WideOr1(WideOr14),
	.av_readdatavalid(av_readdatavalid),
	.out_data_buffer_67(\crosser_003|clock_xer|out_data_buffer[67]~q ),
	.av_readdatavalid1(av_readdatavalid1),
	.av_readdatavalid2(av_readdatavalid2));

usb_system_altera_merlin_slave_translator_7 red_leds_s1_translator(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.reset(altera_reset_synchronizer_int_chain_out),
	.mem_used_1(mem_used_12),
	.always0(always02),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.uav_write(uav_write),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.always1(\router|always1~4_combout ),
	.wait_latency_counter_11(\red_leds_s1_translator|wait_latency_counter[1]~1_combout ),
	.s0_cmd_valid(s0_cmd_valid),
	.read_latency_shift_reg(\red_leds_s1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(\red_leds_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\red_leds_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\red_leds_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\red_leds_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\red_leds_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\red_leds_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\red_leds_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\red_leds_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\red_leds_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\red_leds_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\red_leds_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\red_leds_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\red_leds_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\red_leds_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\red_leds_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\red_leds_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\red_leds_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\red_leds_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_172,readdata_162,readdata_152,readdata_142,readdata_132,readdata_122,readdata_116,readdata_102,readdata_92,readdata_82,readdata_74,readdata_64,readdata_54,readdata_44,readdata_33,readdata_213,readdata_114,readdata_05}),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator all_switches_s1_translator(
	.W_alu_result_7(W_alu_result_7),
	.Equal3(Equal3),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read_latency_shift_reg_0(read_latency_shift_reg_05),
	.uav_write(uav_write),
	.always1(\router|always1~2_combout ),
	.mem_used_1(\all_switches_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\all_switches_s1_translator|wait_latency_counter[1]~1_combout ),
	.waitrequest_reset_override1(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.sink_ready(\cmd_demux|sink_ready~12_combout ),
	.m0_write(\all_switches_s1_agent|m0_write~0_combout ),
	.av_readdata_pre_0(\all_switches_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\all_switches_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\all_switches_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\all_switches_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\all_switches_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\all_switches_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\all_switches_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\all_switches_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\all_switches_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\all_switches_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\all_switches_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\all_switches_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\all_switches_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\all_switches_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\all_switches_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\all_switches_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\all_switches_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\all_switches_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_171,readdata_161,readdata_151,readdata_141,readdata_131,readdata_121,readdata_115,readdata_101,readdata_91,readdata_81,readdata_73,readdata_63,readdata_53,readdata_43,readdata_32,readdata_212,readdata_113,readdata_04}),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator_6 led_s1_translator(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.reset(altera_reset_synchronizer_int_chain_out),
	.mem_used_1(mem_used_11),
	.always0(always01),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.uav_write(uav_write),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.always1(\router|always1~4_combout ),
	.wait_latency_counter_01(\led_s1_translator|wait_latency_counter[0]~1_combout ),
	.s0_cmd_valid(s0_cmd_valid),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(\led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\led_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\led_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\led_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\led_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\led_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\led_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\led_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_71,readdata_61,readdata_51,readdata_41,readdata_34,readdata_210,readdata_110,readdata_02}),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator_5 keycode_s1_translator(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.reset(r_sync_rst),
	.Equal3(Equal3),
	.mem_used_1(mem_used_1),
	.always0(always0),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.read_latency_shift_reg(\keycode_s1_translator|read_latency_shift_reg~2_combout ),
	.sink_in_reset(sink_in_reset),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.read_latency_shift_reg1(\keycode_s1_translator|read_latency_shift_reg~3_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.uav_write(uav_write),
	.s0_cmd_valid(s0_cmd_valid),
	.Equal6(\router|Equal6~2_combout ),
	.av_readdata_pre_0(\keycode_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\keycode_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\keycode_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\keycode_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\keycode_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\keycode_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\keycode_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\keycode_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_72,readdata_62,readdata_52,readdata_42,readdata_35,readdata_211,readdata_112,readdata_03}),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator_2 clocks_pll_slave_translator(
	.reset(r_sync_rst),
	.sink_in_reset(sink_in_reset),
	.read_latency_shift_reg_0(\clocks_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_14),
	.WideOr1(WideOr11),
	.mem(mem1),
	.read_latency_shift_reg(\clocks_pll_slave_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_11,readdata_01}),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator_3 cpu_debug_mem_slave_translator(
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_111,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.sink_in_reset(sink_in_reset),
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_13),
	.local_read(local_read),
	.av_readdata_pre_0(av_readdata_pre_01),
	.av_readdata_pre_1(av_readdata_pre_11),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_11(av_readdata_pre_111),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_30(av_readdata_pre_301),
	.av_readdata_pre_29(av_readdata_pre_29),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator_9 sysid_qsys_0_control_slave_translator(
	.reset(altera_reset_synchronizer_int_chain_out),
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\sysid_qsys_0_control_slave_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ),
	.src_data_68(\cmd_mux_001|src_data[68]~combout ),
	.always1(\router_001|always1~2_combout ),
	.read_latency_shift_reg(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg~1_combout ),
	.WideOr1(\cmd_mux_001|WideOr1~combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata({gnd,\cmd_mux_001|src_data[38]~combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clk(clk_clk));

usb_system_altera_merlin_slave_translator_4 jtag_uart_avalon_jtag_slave_translator(
	.av_readdata_pre_16(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_22(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.reset(r_sync_rst),
	.sink_in_reset(sink_in_reset),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.av_waitrequest(av_waitrequest),
	.sink_ready(sink_ready),
	.av_readdata_pre_0(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,av_readdata_7,av_readdata_6,av_readdata_5,av_readdata_4,av_readdata_3,av_readdata_2,av_readdata_1,av_readdata_0}),
	.av_readdata_pre_9(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_12(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.b_full(b_full),
	.read_0(read_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full1(b_full1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_31(counter_reg_bit_31),
	.counter_reg_bit_21(counter_reg_bit_21),
	.counter_reg_bit_01(counter_reg_bit_01),
	.counter_reg_bit_11(counter_reg_bit_11),
	.counter_reg_bit_41(counter_reg_bit_41),
	.counter_reg_bit_51(counter_reg_bit_51),
	.clk(clk_clk));

usb_system_altera_merlin_master_translator cpu_data_master_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.write_accepted1(write_accepted),
	.sink_in_reset(sink_in_reset),
	.d_read(d_read),
	.read_accepted1(read_accepted),
	.av_ld_getting_data(av_ld_getting_data),
	.uav_write(uav_write),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.WideOr0(\cmd_demux|WideOr0~7_combout ),
	.av_waitrequest(cpu_data_master_waitrequest),
	.s0_cmd_valid(s0_cmd_valid),
	.clk(clk_clk));

usb_system_altera_merlin_master_translator_1 cpu_instruction_master_translator(
	.reset(r_sync_rst),
	.sink_in_reset(sink_in_reset),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_13),
	.mem_used_11(mem_used_14),
	.i_read(i_read),
	.read_accepted1(\cpu_instruction_master_translator|read_accepted~q ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.uav_read(\cpu_instruction_master_translator|uav_read~0_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.Equal2(\router_001|Equal2~2_combout ),
	.saved_grant_11(\cmd_mux_002|saved_grant[1]~q ),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ),
	.av_readdatavalid(av_readdatavalid2),
	.Equal1(\router_001|Equal1~5_combout ),
	.take_in_data(\crosser_001|clock_xer|take_in_data~2_combout ),
	.clk(clk_clk));

usb_system_altera_avalon_sc_fifo all_switches_s1_agent_rsp_fifo(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read_latency_shift_reg_0(read_latency_shift_reg_05),
	.mem_67_0(mem_67_08),
	.mem_used_1(\all_switches_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~13_combout ),
	.clk(clk_clk));

usb_system_altera_merlin_slave_agent all_switches_s1_agent(
	.W_alu_result_7(W_alu_result_7),
	.Equal3(Equal3),
	.always1(\router|always1~2_combout ),
	.mem_used_1(\all_switches_s1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\all_switches_s1_agent|m0_write~0_combout ));

usb_system_altera_avalon_sc_fifo_6 led_s1_agent_rsp_fifo(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.reset(altera_reset_synchronizer_int_chain_out),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.mem_67_0(mem_67_06),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.wait_latency_counter_0(\led_s1_translator|wait_latency_counter[0]~1_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.read_latency_shift_reg(\led_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

usb_system_altera_avalon_sc_fifo_8 sdram_s1_agent_rdata_fifo(
	.clk(wire_pll7_clk_0),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\sdram_s1_agent_rsp_fifo|mem[0][107]~q ),
	.out_valid1(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.WideOr0(\rsp_demux_006|WideOr0~1_combout ),
	.out_payload_0(\sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.out_payload_1(\sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.out_payload_2(\sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.out_payload_3(\sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.out_payload_4(\sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.out_payload_22(\sdram_s1_agent_rdata_fifo|out_payload[22]~q ),
	.out_payload_23(\sdram_s1_agent_rdata_fifo|out_payload[23]~q ),
	.out_payload_24(\sdram_s1_agent_rdata_fifo|out_payload[24]~q ),
	.out_payload_25(\sdram_s1_agent_rdata_fifo|out_payload[25]~q ),
	.out_payload_26(\sdram_s1_agent_rdata_fifo|out_payload[26]~q ),
	.out_payload_11(\sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.out_payload_13(\sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.out_payload_16(\sdram_s1_agent_rdata_fifo|out_payload[16]~q ),
	.out_payload_12(\sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.out_payload_5(\sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.out_payload_14(\sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.out_payload_15(\sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.out_payload_10(\sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.out_payload_9(\sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.out_payload_8(\sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.out_payload_7(\sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.out_payload_6(\sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.out_payload_20(\sdram_s1_agent_rdata_fifo|out_payload[20]~q ),
	.out_payload_18(\sdram_s1_agent_rdata_fifo|out_payload[18]~q ),
	.out_payload_19(\sdram_s1_agent_rdata_fifo|out_payload[19]~q ),
	.out_payload_17(\sdram_s1_agent_rdata_fifo|out_payload[17]~q ),
	.out_payload_21(\sdram_s1_agent_rdata_fifo|out_payload[21]~q ),
	.out_payload_27(\sdram_s1_agent_rdata_fifo|out_payload[27]~q ),
	.out_payload_28(\sdram_s1_agent_rdata_fifo|out_payload[28]~q ),
	.out_payload_31(\sdram_s1_agent_rdata_fifo|out_payload[31]~q ),
	.out_payload_30(\sdram_s1_agent_rdata_fifo|out_payload[30]~q ),
	.out_payload_29(\sdram_s1_agent_rdata_fifo|out_payload[29]~q ),
	.za_valid(za_valid),
	.za_data_0(za_data_0),
	.za_data_1(za_data_1),
	.za_data_2(za_data_2),
	.za_data_3(za_data_3),
	.za_data_4(za_data_4),
	.za_data_22(za_data_22),
	.za_data_23(za_data_23),
	.za_data_24(za_data_24),
	.za_data_25(za_data_25),
	.za_data_26(za_data_26),
	.za_data_11(za_data_11),
	.za_data_13(za_data_13),
	.za_data_16(za_data_16),
	.za_data_12(za_data_12),
	.za_data_5(za_data_5),
	.za_data_14(za_data_14),
	.za_data_15(za_data_15),
	.za_data_10(za_data_10),
	.za_data_9(za_data_9),
	.za_data_8(za_data_8),
	.za_data_7(za_data_7),
	.za_data_6(za_data_6),
	.za_data_20(za_data_20),
	.za_data_18(za_data_18),
	.za_data_19(za_data_19),
	.za_data_17(za_data_17),
	.za_data_21(za_data_21),
	.za_data_27(za_data_27),
	.za_data_28(za_data_28),
	.za_data_31(za_data_31),
	.za_data_30(za_data_30),
	.za_data_29(za_data_29));

usb_system_altera_avalon_sc_fifo_9 sdram_s1_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.last_cycle(last_cycle),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.saved_grant_1(saved_grant_1),
	.WideOr1(WideOr12),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.src_data_68(src_data_68),
	.nonposted_write_endofpacket(\sdram_s1_agent|nonposted_write_endofpacket~0_combout ),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\sdram_s1_agent_rsp_fifo|mem[0][107]~q ),
	.out_valid(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.WideOr0(\rsp_demux_006|WideOr0~1_combout ),
	.mem_67_0(\sdram_s1_agent_rsp_fifo|mem[0][67]~q ),
	.out_data_buffer_86(\crosser_001|clock_xer|out_data_buffer[86]~q ));

usb_system_altera_merlin_slave_agent_8 sdram_s1_agent(
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.WideOr1(WideOr12),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.src_payload(src_payload),
	.src_payload_0(\cmd_mux_006|src_payload[0]~combout ),
	.out_data_buffer_66(\crosser|clock_xer|out_data_buffer[66]~q ),
	.nonposted_write_endofpacket(\sdram_s1_agent|nonposted_write_endofpacket~0_combout ),
	.m0_write(m0_write1));

usb_system_usb_system_mm_interconnect_0_router_001 router_001(
	.F_pc_26(F_pc_26),
	.F_pc_25(F_pc_25),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.Equal1(\router_001|Equal1~4_combout ),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_4(F_pc_4),
	.Equal2(\router_001|Equal2~1_combout ),
	.F_pc_1(F_pc_1),
	.F_pc_3(F_pc_3),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.F_pc_2(F_pc_2),
	.always1(\router_001|always1~1_combout ),
	.Equal21(\router_001|Equal2~2_combout ),
	.always11(\router_001|always1~2_combout ),
	.Equal11(\router_001|Equal1~5_combout ));

usb_system_usb_system_mm_interconnect_0_router router(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_3(W_alu_result_3),
	.Equal1(\router|Equal1~0_combout ),
	.Equal3(Equal3),
	.Equal6(Equal6),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.Equal2(\router|Equal2~5_combout ),
	.always1(\router|always1~2_combout ),
	.Equal11(\router|Equal1~2_combout ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.always11(\router|always1~3_combout ),
	.Equal9(\router|Equal9~0_combout ),
	.Equal91(Equal9),
	.always12(\router|always1~4_combout ),
	.Equal5(\router|Equal5~0_combout ),
	.Equal31(\router|Equal3~6_combout ),
	.Equal7(\router|Equal7~0_combout ),
	.Equal61(\router|Equal6~2_combout ),
	.always13(\router|always1~5_combout ),
	.Equal12(\router|Equal1~3_combout ),
	.always14(\router|always1~6_combout ));

usb_system_altera_avalon_sc_fifo_7 red_leds_s1_agent_rsp_fifo(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.reset(altera_reset_synchronizer_int_chain_out),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_67_0(mem_67_07),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.wait_latency_counter_1(\red_leds_s1_translator|wait_latency_counter[1]~1_combout ),
	.Equal3(\router|Equal3~6_combout ),
	.read_latency_shift_reg(\red_leds_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

usb_system_altera_avalon_st_handshake_clock_crosser_3 crosser_003(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.out_data_toggle_flopped(\crosser_003|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_003|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(out_valid2),
	.out_data_buffer_67(\crosser_003|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(\crosser_003|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(out_data_buffer_4),
	.in_data_toggle(\crosser_003|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_003|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.always0(\router_008|always0~0_combout ),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(\crosser_003|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_20(\crosser_003|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_21(\crosser_003|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.mem_67_0(\sdram_s1_agent_rsp_fifo|mem[0][67]~q ),
	.take_in_data(\crosser_002|clock_xer|take_in_data~0_combout ),
	.out_payload_0(\sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.out_payload_1(\sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.out_payload_2(\sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.out_payload_3(\sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.out_payload_4(\sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.out_payload_22(\sdram_s1_agent_rdata_fifo|out_payload[22]~q ),
	.out_payload_23(\sdram_s1_agent_rdata_fifo|out_payload[23]~q ),
	.out_payload_24(\sdram_s1_agent_rdata_fifo|out_payload[24]~q ),
	.out_payload_25(\sdram_s1_agent_rdata_fifo|out_payload[25]~q ),
	.out_payload_26(\sdram_s1_agent_rdata_fifo|out_payload[26]~q ),
	.out_payload_11(\sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.out_payload_13(\sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.out_payload_16(\sdram_s1_agent_rdata_fifo|out_payload[16]~q ),
	.out_payload_12(\sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.out_payload_5(\sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.out_payload_14(\sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.out_payload_15(\sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.out_payload_10(\sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.out_payload_9(\sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.out_payload_8(\sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.out_payload_7(\sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.out_payload_6(\sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.out_payload_20(\sdram_s1_agent_rdata_fifo|out_payload[20]~q ),
	.out_payload_18(\sdram_s1_agent_rdata_fifo|out_payload[18]~q ),
	.out_payload_19(\sdram_s1_agent_rdata_fifo|out_payload[19]~q ),
	.out_payload_17(\sdram_s1_agent_rdata_fifo|out_payload[17]~q ),
	.out_payload_21(\sdram_s1_agent_rdata_fifo|out_payload[21]~q ),
	.out_payload_27(\sdram_s1_agent_rdata_fifo|out_payload[27]~q ),
	.out_payload_28(\sdram_s1_agent_rdata_fifo|out_payload[28]~q ),
	.out_payload_31(\sdram_s1_agent_rdata_fifo|out_payload[31]~q ),
	.out_payload_30(\sdram_s1_agent_rdata_fifo|out_payload[30]~q ),
	.out_payload_29(\sdram_s1_agent_rdata_fifo|out_payload[29]~q ),
	.clk_clk(clk_clk));

usb_system_altera_avalon_st_handshake_clock_crosser_2 crosser_002(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.out_data_toggle_flopped(\crosser_002|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_002|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(out_valid1),
	.out_data_buffer_67(out_data_buffer_67),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\sdram_s1_agent_rsp_fifo|mem[0][107]~q ),
	.out_valid1(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.in_data_toggle(\crosser_002|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_002|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.always0(\router_008|always0~0_combout ),
	.out_data_buffer_0(\crosser_002|clock_xer|out_data_buffer[0]~q ),
	.mem_67_0(\sdram_s1_agent_rsp_fifo|mem[0][67]~q ),
	.take_in_data(\crosser_002|clock_xer|take_in_data~0_combout ),
	.out_data_buffer_1(\crosser_002|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser_002|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser_002|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser_002|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser_002|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser_002|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser_002|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_8(\crosser_002|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_9(\crosser_002|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_10(\crosser_002|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_11(\crosser_002|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_12(\crosser_002|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_13(\crosser_002|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_14(\crosser_002|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_15(\crosser_002|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_16(\crosser_002|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_17(\crosser_002|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_18(\crosser_002|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_23(\crosser_002|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_22(\crosser_002|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_21(\crosser_002|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_20(\crosser_002|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_19(\crosser_002|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_24(out_data_buffer_241),
	.out_data_buffer_28(out_data_buffer_281),
	.out_data_buffer_27(out_data_buffer_271),
	.out_data_buffer_26(out_data_buffer_261),
	.out_data_buffer_25(out_data_buffer_251),
	.out_payload_0(\sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.out_payload_1(\sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.out_payload_2(\sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.out_payload_3(\sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.out_payload_4(\sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.out_payload_22(\sdram_s1_agent_rdata_fifo|out_payload[22]~q ),
	.out_payload_23(\sdram_s1_agent_rdata_fifo|out_payload[23]~q ),
	.out_payload_24(\sdram_s1_agent_rdata_fifo|out_payload[24]~q ),
	.out_payload_25(\sdram_s1_agent_rdata_fifo|out_payload[25]~q ),
	.out_payload_26(\sdram_s1_agent_rdata_fifo|out_payload[26]~q ),
	.out_payload_11(\sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.out_payload_13(\sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.out_payload_16(\sdram_s1_agent_rdata_fifo|out_payload[16]~q ),
	.out_payload_12(\sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.out_payload_5(\sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.out_payload_14(\sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.out_payload_15(\sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.out_payload_10(\sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.out_payload_9(\sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.out_payload_8(\sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.out_payload_7(\sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.out_payload_6(\sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.out_payload_20(\sdram_s1_agent_rdata_fifo|out_payload[20]~q ),
	.out_payload_18(\sdram_s1_agent_rdata_fifo|out_payload[18]~q ),
	.out_payload_19(\sdram_s1_agent_rdata_fifo|out_payload[19]~q ),
	.out_payload_17(\sdram_s1_agent_rdata_fifo|out_payload[17]~q ),
	.out_payload_21(\sdram_s1_agent_rdata_fifo|out_payload[21]~q ),
	.out_data_buffer_31(out_data_buffer_311),
	.out_payload_27(\sdram_s1_agent_rdata_fifo|out_payload[27]~q ),
	.out_data_buffer_30(out_data_buffer_301),
	.out_data_buffer_29(out_data_buffer_291),
	.out_payload_28(\sdram_s1_agent_rdata_fifo|out_payload[28]~q ),
	.out_payload_31(\sdram_s1_agent_rdata_fifo|out_payload[31]~q ),
	.out_payload_30(\sdram_s1_agent_rdata_fifo|out_payload[30]~q ),
	.out_payload_29(\sdram_s1_agent_rdata_fifo|out_payload[29]~q ),
	.clk_clk(clk_clk));

usb_system_altera_avalon_st_handshake_clock_crosser_1 crosser_001(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_4(F_pc_4),
	.F_pc_1(F_pc_1),
	.F_pc_3(F_pc_3),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.F_pc_2(F_pc_2),
	.Equal2(\router_001|Equal2~2_combout ),
	.F_pc_0(F_pc_0),
	.last_cycle(last_cycle),
	.saved_grant_1(saved_grant_1),
	.out_valid(\crosser_001|clock_xer|out_valid~combout ),
	.out_data_buffer_68(\crosser_001|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_48(\crosser_001|clock_xer|out_data_buffer[48]~q ),
	.out_data_buffer_62(\crosser_001|clock_xer|out_data_buffer[62]~q ),
	.out_data_buffer_49(\crosser_001|clock_xer|out_data_buffer[49]~q ),
	.out_data_buffer_51(\crosser_001|clock_xer|out_data_buffer[51]~q ),
	.out_data_buffer_50(\crosser_001|clock_xer|out_data_buffer[50]~q ),
	.out_data_buffer_53(\crosser_001|clock_xer|out_data_buffer[53]~q ),
	.out_data_buffer_52(\crosser_001|clock_xer|out_data_buffer[52]~q ),
	.out_data_buffer_55(\crosser_001|clock_xer|out_data_buffer[55]~q ),
	.out_data_buffer_54(\crosser_001|clock_xer|out_data_buffer[54]~q ),
	.out_data_buffer_57(\crosser_001|clock_xer|out_data_buffer[57]~q ),
	.out_data_buffer_56(\crosser_001|clock_xer|out_data_buffer[56]~q ),
	.out_data_buffer_59(\crosser_001|clock_xer|out_data_buffer[59]~q ),
	.out_data_buffer_58(\crosser_001|clock_xer|out_data_buffer[58]~q ),
	.out_data_buffer_61(\crosser_001|clock_xer|out_data_buffer[61]~q ),
	.out_data_buffer_60(\crosser_001|clock_xer|out_data_buffer[60]~q ),
	.out_data_buffer_38(\crosser_001|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser_001|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_40(\crosser_001|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_41(\crosser_001|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_42(\crosser_001|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_43(\crosser_001|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_44(\crosser_001|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_45(\crosser_001|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_46(\crosser_001|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_47(\crosser_001|clock_xer|out_data_buffer[47]~q ),
	.out_data_buffer_32(out_data_buffer_321),
	.out_data_buffer_33(out_data_buffer_331),
	.out_data_buffer_34(out_data_buffer_341),
	.out_data_buffer_35(out_data_buffer_351),
	.always1(\router_001|always1~2_combout ),
	.Equal1(\router_001|Equal1~5_combout ),
	.take_in_data(\crosser_001|clock_xer|take_in_data~2_combout ),
	.out_data_buffer_107(\crosser_001|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_86(\crosser_001|clock_xer|out_data_buffer[86]~q ),
	.clk_clk(clk_clk));

usb_system_altera_avalon_st_handshake_clock_crosser crosser(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.uav_write(uav_write),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.sink_ready(\cmd_demux|sink_ready~7_combout ),
	.in_data_toggle(\crosser|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.s0_cmd_valid(s0_cmd_valid),
	.last_cycle(last_cycle),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.out_data_toggle_flopped(\crosser|clock_xer|out_data_toggle_flopped~q ),
	.dreg_01(\crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(\crosser|clock_xer|out_valid~combout ),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_68(\crosser|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_48(\crosser|clock_xer|out_data_buffer[48]~q ),
	.out_data_buffer_62(\crosser|clock_xer|out_data_buffer[62]~q ),
	.out_data_buffer_49(\crosser|clock_xer|out_data_buffer[49]~q ),
	.out_data_buffer_51(\crosser|clock_xer|out_data_buffer[51]~q ),
	.out_data_buffer_50(\crosser|clock_xer|out_data_buffer[50]~q ),
	.out_data_buffer_53(\crosser|clock_xer|out_data_buffer[53]~q ),
	.out_data_buffer_52(\crosser|clock_xer|out_data_buffer[52]~q ),
	.out_data_buffer_55(\crosser|clock_xer|out_data_buffer[55]~q ),
	.out_data_buffer_54(\crosser|clock_xer|out_data_buffer[54]~q ),
	.out_data_buffer_57(\crosser|clock_xer|out_data_buffer[57]~q ),
	.out_data_buffer_56(\crosser|clock_xer|out_data_buffer[56]~q ),
	.out_data_buffer_59(\crosser|clock_xer|out_data_buffer[59]~q ),
	.out_data_buffer_58(\crosser|clock_xer|out_data_buffer[58]~q ),
	.out_data_buffer_61(\crosser|clock_xer|out_data_buffer[61]~q ),
	.out_data_buffer_60(\crosser|clock_xer|out_data_buffer[60]~q ),
	.out_data_buffer_38(\crosser|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_40(\crosser|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_41(\crosser|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_42(\crosser|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_43(\crosser|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_44(\crosser|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_45(\crosser|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_46(\crosser|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_47(\crosser|clock_xer|out_data_buffer[47]~q ),
	.out_data_buffer_32(out_data_buffer_32),
	.out_data_buffer_33(out_data_buffer_33),
	.out_data_buffer_34(out_data_buffer_34),
	.out_data_buffer_35(out_data_buffer_35),
	.sink_ready1(\cmd_demux|sink_ready~14_combout ),
	.out_data_buffer_107(\crosser|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_66(\crosser|clock_xer|out_data_buffer[66]~q ),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.out_data_buffer_0(\crosser|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_8(\crosser|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_9(\crosser|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_10(\crosser|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_11(\crosser|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_12(\crosser|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_13(\crosser|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_14(\crosser|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_15(\crosser|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_16(\crosser|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_17(\crosser|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_18(\crosser|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_19(\crosser|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_20(\crosser|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_21(\crosser|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_22(\crosser|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_23(\crosser|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_24(\crosser|clock_xer|out_data_buffer[24]~q ),
	.out_data_buffer_25(\crosser|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_26(\crosser|clock_xer|out_data_buffer[26]~q ),
	.out_data_buffer_27(\crosser|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_28(\crosser|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_29(\crosser|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_30(\crosser|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_31(\crosser|clock_xer|out_data_buffer[31]~q ),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.clk_clk(clk_clk));

usb_system_usb_system_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.read_latency_shift_reg_01(\clocks_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_01(\clocks_pll_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_01(\clocks_pll_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src1_valid(src1_valid),
	.src_payload(src_payload1),
	.out_data_toggle_flopped(\crosser_003|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_003|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(out_valid2),
	.src_payload1(src_payload2),
	.WideOr1(WideOr14),
	.out_data_buffer_3(\crosser_003|clock_xer|out_data_buffer[3]~q ),
	.src_payload2(src_payload3),
	.out_data_buffer_16(\crosser_003|clock_xer|out_data_buffer[16]~q ),
	.src_payload3(src_payload4),
	.out_data_buffer_20(\crosser_003|clock_xer|out_data_buffer[20]~q ),
	.src_payload4(src_payload5),
	.out_data_buffer_21(\crosser_003|clock_xer|out_data_buffer[21]~q ),
	.src_payload5(src_payload6));

usb_system_usb_system_mm_interconnect_0_rsp_mux rsp_mux(
	.av_readdata_pre_16(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_22(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.out_valid(out_valid),
	.read_latency_shift_reg_02(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid),
	.read_latency_shift_reg_03(read_latency_shift_reg_02),
	.read_latency_shift_reg_04(read_latency_shift_reg_03),
	.mem_86_01(mem_86_0),
	.mem_68_01(mem_68_0),
	.src0_valid1(src0_valid1),
	.read_latency_shift_reg_05(\clocks_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_02(\clocks_pll_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_02(\clocks_pll_slave_agent_rsp_fifo|mem[0][68]~q ),
	.read_latency_shift_reg_06(read_latency_shift_reg_04),
	.read_latency_shift_reg_07(read_latency_shift_reg_05),
	.out_data_toggle_flopped(\crosser_002|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_002|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.WideOr11(WideOr1),
	.src0_valid2(src0_valid2),
	.out_valid1(out_valid1),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_01(av_readdata_pre_01),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_02(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.out_payload_0(out_payload_0),
	.av_readdata_pre_03(\led_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_04(\keycode_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_05(\all_switches_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_06(\red_leds_s1_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_0(\crosser_002|clock_xer|out_data_buffer[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_221(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_111(av_readdata_pre_111),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_161(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_201(av_readdata_pre_20),
	.av_readdata_pre_181(av_readdata_pre_18),
	.av_readdata_pre_191(av_readdata_pre_19),
	.av_readdata_pre_171(av_readdata_pre_17),
	.av_readdata_pre_211(av_readdata_pre_21),
	.av_readdata_pre_110(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.out_payload_1(out_payload_1),
	.av_readdata_pre_112(\led_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_113(\keycode_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_114(\all_switches_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_115(\red_leds_s1_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_1(\crosser_002|clock_xer|out_data_buffer[1]~q ),
	.src_data_1(src_data_1),
	.src_payload(src_payload7),
	.av_readdata_pre_24(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.out_payload_2(out_payload_2),
	.av_readdata_pre_25(\led_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_26(\keycode_s1_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_27(\all_switches_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_28(\red_leds_s1_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_2(\crosser_002|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_31(\all_switches_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\red_leds_s1_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_33(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.out_payload_3(out_payload_3),
	.av_readdata_pre_34(\led_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_35(\keycode_s1_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_3(\crosser_002|clock_xer|out_data_buffer[3]~q ),
	.src_data_31(src_data_31),
	.av_readdata_pre_41(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.out_payload_4(out_payload_4),
	.av_readdata_pre_42(\led_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\keycode_s1_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_44(\all_switches_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_45(\red_leds_s1_translator|av_readdata_pre[4]~q ),
	.out_data_buffer_4(\crosser_002|clock_xer|out_data_buffer[4]~q ),
	.av_readdata_pre_51(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.out_payload_5(out_payload_5),
	.av_readdata_pre_52(\led_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\keycode_s1_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_54(\all_switches_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_55(\red_leds_s1_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_5(\crosser_002|clock_xer|out_data_buffer[5]~q ),
	.av_readdata_pre_61(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.out_payload_6(out_payload_6),
	.av_readdata_pre_62(\led_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\keycode_s1_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_64(\all_switches_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_65(\red_leds_s1_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_6(\crosser_002|clock_xer|out_data_buffer[6]~q ),
	.av_readdata_pre_71(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.out_payload_7(out_payload_7),
	.av_readdata_pre_72(\led_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\keycode_s1_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_74(\all_switches_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_75(\red_leds_s1_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_7(\crosser_002|clock_xer|out_data_buffer[7]~q ),
	.av_readdata_pre_81(\all_switches_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\red_leds_s1_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_8(\crosser_002|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_83(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.out_payload_8(out_payload_8),
	.src_data_8(src_data_8),
	.av_readdata_pre_91(\all_switches_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\red_leds_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_93(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.out_payload_9(out_payload_9),
	.out_data_buffer_9(\crosser_002|clock_xer|out_data_buffer[9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_101(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.out_payload_10(out_payload_10),
	.av_readdata_pre_102(\all_switches_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_103(\red_leds_s1_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_10(\crosser_002|clock_xer|out_data_buffer[10]~q ),
	.src_data_10(src_data_10),
	.av_readdata_pre_116(\all_switches_s1_translator|av_readdata_pre[11]~q ),
	.out_payload_11(out_payload_11),
	.out_data_buffer_11(\crosser_002|clock_xer|out_data_buffer[11]~q ),
	.av_readdata_pre_117(\red_leds_s1_translator|av_readdata_pre[11]~q ),
	.src_data_11(src_data_11),
	.av_readdata_pre_121(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.out_payload_12(out_payload_12),
	.av_readdata_pre_122(\all_switches_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_123(\red_leds_s1_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\crosser_002|clock_xer|out_data_buffer[12]~q ),
	.src_data_12(src_data_12),
	.av_readdata_pre_131(\all_switches_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_132(\red_leds_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_133(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.out_payload_13(out_payload_13),
	.out_data_buffer_13(\crosser_002|clock_xer|out_data_buffer[13]~q ),
	.src_data_13(src_data_13),
	.av_readdata_pre_141(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.out_payload_14(out_payload_14),
	.av_readdata_pre_142(\all_switches_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_143(\red_leds_s1_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_14(\crosser_002|clock_xer|out_data_buffer[14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_151(\all_switches_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_152(\red_leds_s1_translator|av_readdata_pre[15]~q ),
	.out_data_buffer_15(\crosser_002|clock_xer|out_data_buffer[15]~q ),
	.av_readdata_pre_153(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.out_payload_15(out_payload_15),
	.src_data_15(src_data_15),
	.av_readdata_pre_162(\all_switches_s1_translator|av_readdata_pre[16]~q ),
	.out_data_buffer_16(\crosser_002|clock_xer|out_data_buffer[16]~q ),
	.av_readdata_pre_163(\red_leds_s1_translator|av_readdata_pre[16]~q ),
	.src_data_16(src_data_16),
	.av_readdata_pre_172(\all_switches_s1_translator|av_readdata_pre[17]~q ),
	.out_data_buffer_17(\crosser_002|clock_xer|out_data_buffer[17]~q ),
	.av_readdata_pre_173(\red_leds_s1_translator|av_readdata_pre[17]~q ),
	.src_data_17(src_data_17),
	.out_data_buffer_18(\crosser_002|clock_xer|out_data_buffer[18]~q ),
	.src_payload1(src_payload40),
	.out_data_buffer_23(\crosser_002|clock_xer|out_data_buffer[23]~q ),
	.src_payload2(src_payload41),
	.out_data_buffer_22(\crosser_002|clock_xer|out_data_buffer[22]~q ),
	.src_payload3(src_payload42),
	.out_data_buffer_21(\crosser_002|clock_xer|out_data_buffer[21]~q ),
	.src_payload4(src_payload43),
	.out_data_buffer_20(\crosser_002|clock_xer|out_data_buffer[20]~q ),
	.src_payload5(src_payload44),
	.out_data_buffer_19(\crosser_002|clock_xer|out_data_buffer[19]~q ),
	.src_payload6(src_payload45),
	.src_data_21(src_data_21),
	.src_data_41(src_data_410),
	.src_data_51(src_data_510),
	.src_data_61(src_data_63),
	.src_data_71(src_data_71));

usb_system_usb_system_mm_interconnect_0_rsp_demux_001_3 rsp_demux_006(
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.in_data_toggle(\crosser_003|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_003|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.in_data_toggle1(\crosser_002|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_002|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.always0(\router_008|always0~0_combout ),
	.WideOr0(\rsp_demux_006|WideOr0~1_combout ));

usb_system_usb_system_mm_interconnect_0_rsp_demux_001_2 rsp_demux_003(
	.read_latency_shift_reg_0(\clocks_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\clocks_pll_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\clocks_pll_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid2));

usb_system_usb_system_mm_interconnect_0_rsp_demux_001_1 rsp_demux_002(
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid));

usb_system_usb_system_mm_interconnect_0_rsp_demux_001 rsp_demux_001(
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid));

usb_system_usb_system_mm_interconnect_0_cmd_mux_001_3 cmd_mux_006(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.last_cycle(last_cycle),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.saved_grant_1(saved_grant_1),
	.out_valid(\crosser_001|clock_xer|out_valid~combout ),
	.out_data_toggle_flopped(\crosser|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid1(\crosser|clock_xer|out_valid~combout ),
	.WideOr11(WideOr12),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.src_payload(src_payload),
	.out_data_buffer_68(\crosser_001|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_681(\crosser|clock_xer|out_data_buffer[68]~q ),
	.src_data_68(src_data_68),
	.out_data_buffer_48(\crosser_001|clock_xer|out_data_buffer[48]~q ),
	.out_data_buffer_481(\crosser|clock_xer|out_data_buffer[48]~q ),
	.src_data_48(src_data_48),
	.out_data_buffer_62(\crosser_001|clock_xer|out_data_buffer[62]~q ),
	.out_data_buffer_621(\crosser|clock_xer|out_data_buffer[62]~q ),
	.src_data_62(src_data_62),
	.out_data_buffer_49(\crosser_001|clock_xer|out_data_buffer[49]~q ),
	.out_data_buffer_491(\crosser|clock_xer|out_data_buffer[49]~q ),
	.src_data_49(src_data_49),
	.out_data_buffer_51(\crosser_001|clock_xer|out_data_buffer[51]~q ),
	.out_data_buffer_511(\crosser|clock_xer|out_data_buffer[51]~q ),
	.src_data_51(src_data_51),
	.out_data_buffer_50(\crosser_001|clock_xer|out_data_buffer[50]~q ),
	.out_data_buffer_501(\crosser|clock_xer|out_data_buffer[50]~q ),
	.src_data_50(src_data_50),
	.out_data_buffer_53(\crosser_001|clock_xer|out_data_buffer[53]~q ),
	.out_data_buffer_531(\crosser|clock_xer|out_data_buffer[53]~q ),
	.src_data_53(src_data_53),
	.out_data_buffer_52(\crosser_001|clock_xer|out_data_buffer[52]~q ),
	.out_data_buffer_521(\crosser|clock_xer|out_data_buffer[52]~q ),
	.src_data_52(src_data_52),
	.out_data_buffer_55(\crosser_001|clock_xer|out_data_buffer[55]~q ),
	.out_data_buffer_551(\crosser|clock_xer|out_data_buffer[55]~q ),
	.src_data_55(src_data_55),
	.out_data_buffer_54(\crosser_001|clock_xer|out_data_buffer[54]~q ),
	.out_data_buffer_541(\crosser|clock_xer|out_data_buffer[54]~q ),
	.src_data_54(src_data_54),
	.out_data_buffer_57(\crosser_001|clock_xer|out_data_buffer[57]~q ),
	.out_data_buffer_571(\crosser|clock_xer|out_data_buffer[57]~q ),
	.src_data_57(src_data_57),
	.out_data_buffer_56(\crosser_001|clock_xer|out_data_buffer[56]~q ),
	.out_data_buffer_561(\crosser|clock_xer|out_data_buffer[56]~q ),
	.src_data_56(src_data_56),
	.out_data_buffer_59(\crosser_001|clock_xer|out_data_buffer[59]~q ),
	.out_data_buffer_591(\crosser|clock_xer|out_data_buffer[59]~q ),
	.src_data_59(src_data_59),
	.out_data_buffer_58(\crosser_001|clock_xer|out_data_buffer[58]~q ),
	.out_data_buffer_581(\crosser|clock_xer|out_data_buffer[58]~q ),
	.src_data_58(src_data_58),
	.out_data_buffer_61(\crosser_001|clock_xer|out_data_buffer[61]~q ),
	.out_data_buffer_611(\crosser|clock_xer|out_data_buffer[61]~q ),
	.src_data_61(src_data_61),
	.out_data_buffer_60(\crosser_001|clock_xer|out_data_buffer[60]~q ),
	.out_data_buffer_601(\crosser|clock_xer|out_data_buffer[60]~q ),
	.src_data_60(src_data_60),
	.out_data_buffer_38(\crosser_001|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_381(\crosser|clock_xer|out_data_buffer[38]~q ),
	.src_data_38(src_data_381),
	.out_data_buffer_39(\crosser_001|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_391(\crosser|clock_xer|out_data_buffer[39]~q ),
	.src_data_39(src_data_391),
	.out_data_buffer_40(\crosser_001|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_401(\crosser|clock_xer|out_data_buffer[40]~q ),
	.src_data_40(src_data_40),
	.out_data_buffer_41(\crosser_001|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_411(\crosser|clock_xer|out_data_buffer[41]~q ),
	.src_data_41(src_data_41),
	.out_data_buffer_42(\crosser_001|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_421(\crosser|clock_xer|out_data_buffer[42]~q ),
	.src_data_42(src_data_42),
	.out_data_buffer_43(\crosser_001|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_431(\crosser|clock_xer|out_data_buffer[43]~q ),
	.src_data_43(src_data_43),
	.out_data_buffer_44(\crosser_001|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_441(\crosser|clock_xer|out_data_buffer[44]~q ),
	.src_data_44(src_data_44),
	.out_data_buffer_45(\crosser_001|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_451(\crosser|clock_xer|out_data_buffer[45]~q ),
	.src_data_45(src_data_45),
	.out_data_buffer_46(\crosser_001|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_461(\crosser|clock_xer|out_data_buffer[46]~q ),
	.src_data_46(src_data_46),
	.out_data_buffer_47(\crosser_001|clock_xer|out_data_buffer[47]~q ),
	.out_data_buffer_471(\crosser|clock_xer|out_data_buffer[47]~q ),
	.src_data_47(src_data_47),
	.out_data_buffer_107(\crosser_001|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_1071(\crosser|clock_xer|out_data_buffer[107]~q ),
	.src_payload_0(\cmd_mux_006|src_payload[0]~combout ),
	.out_data_buffer_0(\crosser|clock_xer|out_data_buffer[0]~q ),
	.src_payload1(src_payload8),
	.out_data_buffer_1(\crosser|clock_xer|out_data_buffer[1]~q ),
	.src_payload2(src_payload9),
	.out_data_buffer_2(\crosser|clock_xer|out_data_buffer[2]~q ),
	.src_payload3(src_payload10),
	.out_data_buffer_3(\crosser|clock_xer|out_data_buffer[3]~q ),
	.src_payload4(src_payload11),
	.out_data_buffer_4(\crosser|clock_xer|out_data_buffer[4]~q ),
	.src_payload5(src_payload12),
	.out_data_buffer_5(\crosser|clock_xer|out_data_buffer[5]~q ),
	.src_payload6(src_payload13),
	.out_data_buffer_6(\crosser|clock_xer|out_data_buffer[6]~q ),
	.src_payload7(src_payload14),
	.out_data_buffer_7(\crosser|clock_xer|out_data_buffer[7]~q ),
	.src_payload8(src_payload15),
	.out_data_buffer_8(\crosser|clock_xer|out_data_buffer[8]~q ),
	.src_payload9(src_payload16),
	.out_data_buffer_9(\crosser|clock_xer|out_data_buffer[9]~q ),
	.src_payload10(src_payload17),
	.out_data_buffer_10(\crosser|clock_xer|out_data_buffer[10]~q ),
	.src_payload11(src_payload18),
	.out_data_buffer_11(\crosser|clock_xer|out_data_buffer[11]~q ),
	.src_payload12(src_payload19),
	.out_data_buffer_12(\crosser|clock_xer|out_data_buffer[12]~q ),
	.src_payload13(src_payload20),
	.out_data_buffer_13(\crosser|clock_xer|out_data_buffer[13]~q ),
	.src_payload14(src_payload21),
	.out_data_buffer_14(\crosser|clock_xer|out_data_buffer[14]~q ),
	.src_payload15(src_payload22),
	.out_data_buffer_15(\crosser|clock_xer|out_data_buffer[15]~q ),
	.src_payload16(src_payload23),
	.out_data_buffer_16(\crosser|clock_xer|out_data_buffer[16]~q ),
	.src_payload17(src_payload24),
	.out_data_buffer_17(\crosser|clock_xer|out_data_buffer[17]~q ),
	.src_payload18(src_payload25),
	.out_data_buffer_18(\crosser|clock_xer|out_data_buffer[18]~q ),
	.src_payload19(src_payload26),
	.out_data_buffer_19(\crosser|clock_xer|out_data_buffer[19]~q ),
	.src_payload20(src_payload27),
	.out_data_buffer_20(\crosser|clock_xer|out_data_buffer[20]~q ),
	.src_payload21(src_payload28),
	.out_data_buffer_21(\crosser|clock_xer|out_data_buffer[21]~q ),
	.src_payload22(src_payload29),
	.out_data_buffer_22(\crosser|clock_xer|out_data_buffer[22]~q ),
	.src_payload23(src_payload30),
	.out_data_buffer_23(\crosser|clock_xer|out_data_buffer[23]~q ),
	.src_payload24(src_payload31),
	.out_data_buffer_24(\crosser|clock_xer|out_data_buffer[24]~q ),
	.src_payload25(src_payload32),
	.out_data_buffer_25(\crosser|clock_xer|out_data_buffer[25]~q ),
	.src_payload26(src_payload33),
	.out_data_buffer_26(\crosser|clock_xer|out_data_buffer[26]~q ),
	.src_payload27(src_payload34),
	.out_data_buffer_27(\crosser|clock_xer|out_data_buffer[27]~q ),
	.src_payload28(src_payload35),
	.out_data_buffer_28(\crosser|clock_xer|out_data_buffer[28]~q ),
	.src_payload29(src_payload36),
	.out_data_buffer_29(\crosser|clock_xer|out_data_buffer[29]~q ),
	.src_payload30(src_payload37),
	.out_data_buffer_30(\crosser|clock_xer|out_data_buffer[30]~q ),
	.src_payload31(src_payload38),
	.out_data_buffer_31(\crosser|clock_xer|out_data_buffer[31]~q ),
	.src_payload32(src_payload39));

usb_system_usb_system_mm_interconnect_0_cmd_mux_001_2 cmd_mux_003(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.r_sync_rst(r_sync_rst),
	.Equal6(Equal6),
	.sink_in_reset(sink_in_reset),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(mem_used_14),
	.F_pc_1(F_pc_1),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.s0_cmd_valid(s0_cmd_valid),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.Equal2(\router_001|Equal2~2_combout ),
	.Equal7(\router|Equal7~0_combout ),
	.WideOr11(WideOr11),
	.F_pc_0(F_pc_0),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ),
	.clk_clk(clk_clk));

usb_system_usb_system_mm_interconnect_0_cmd_mux_001_1 cmd_mux_002(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.Equal2(\router|Equal2~5_combout ),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_13),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_5(F_pc_5),
	.F_pc_6(F_pc_6),
	.F_pc_4(F_pc_4),
	.F_pc_1(F_pc_1),
	.F_pc_3(F_pc_3),
	.F_pc_2(F_pc_2),
	.s0_cmd_valid(s0_cmd_valid),
	.F_pc_0(F_pc_0),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.WideOr11(WideOr13),
	.hbreak_enabled(hbreak_enabled),
	.src_data_46(src_data_461),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.src_payload(src_payload46),
	.src_payload1(src_payload47),
	.src_data_38(src_data_382),
	.src_data_39(src_data_392),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_32(src_data_32),
	.src_payload2(src_payload48),
	.src_payload3(src_payload49),
	.src_payload4(src_payload50),
	.src_payload5(src_payload51),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.src_payload6(src_payload52),
	.src_payload7(src_payload53),
	.src_payload8(src_payload54),
	.src_data_34(src_data_34),
	.src_payload9(src_payload55),
	.src_payload10(src_payload56),
	.src_payload11(src_payload57),
	.src_data_35(src_data_35),
	.src_payload12(src_payload58),
	.src_payload13(src_payload59),
	.src_payload14(src_payload60),
	.src_data_33(src_data_33),
	.src_payload15(src_payload61),
	.src_payload16(src_payload62),
	.src_payload17(src_payload63),
	.src_payload18(src_payload64),
	.src_payload19(src_payload65),
	.src_payload20(src_payload66),
	.src_payload21(src_payload67),
	.src_payload22(src_payload68),
	.src_payload23(src_payload69),
	.src_payload24(src_payload70),
	.src_payload25(src_payload71),
	.src_payload26(src_payload72),
	.src_payload27(src_payload73),
	.src_payload28(src_payload74),
	.src_payload29(src_payload75),
	.src_payload30(src_payload76),
	.src_payload31(src_payload77),
	.src_payload32(src_payload78),
	.clk_clk(clk_clk));

usb_system_usb_system_mm_interconnect_0_cmd_mux_001 cmd_mux_001(
	.W_alu_result_2(W_alu_result_2),
	.Equal6(Equal6),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.uav_read(\cpu_data_master_translator|uav_read~0_combout ),
	.always1(\router|always1~3_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.Equal1(\router_001|Equal1~4_combout ),
	.Equal2(\router_001|Equal2~1_combout ),
	.always11(\router_001|always1~1_combout ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.uav_read1(\cpu_instruction_master_translator|uav_read~0_combout ),
	.F_pc_0(F_pc_0),
	.src_data_68(\cmd_mux_001|src_data[68]~combout ),
	.always12(\router_001|always1~2_combout ),
	.always13(\router|always1~6_combout ),
	.WideOr11(\cmd_mux_001|WideOr1~combout ),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_data_38(\cmd_mux_001|src_data[38]~combout ),
	.clk_clk(clk_clk));

usb_system_usb_system_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.Equal1(\router_001|Equal1~4_combout ),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.i_read(i_read),
	.read_accepted(\cpu_instruction_master_translator|read_accepted~q ),
	.uav_read(\cpu_instruction_master_translator|uav_read~0_combout ),
	.Equal2(\router_001|Equal2~2_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ));

usb_system_usb_system_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_5(W_alu_result_5),
	.Equal3(Equal3),
	.mem_used_1(mem_used_1),
	.always0(always01),
	.always01(always02),
	.read_latency_shift_reg(\keycode_s1_translator|read_latency_shift_reg~2_combout ),
	.sink_in_reset(sink_in_reset),
	.Equal2(\router|Equal2~5_combout ),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(waitrequest),
	.mem_used_11(mem_used_13),
	.always1(\router|always1~2_combout ),
	.mem_used_12(\all_switches_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\all_switches_s1_translator|wait_latency_counter[1]~1_combout ),
	.waitrequest_reset_override(\all_switches_s1_translator|waitrequest_reset_override~q ),
	.saved_grant_01(\cmd_mux_003|saved_grant[0]~q ),
	.mem_used_13(mem_used_14),
	.full(full),
	.mem_used_128(\clock_crossing_io_s0_agent_rsp_fifo|mem_used[128]~q ),
	.Equal1(\router|Equal1~2_combout ),
	.saved_grant_02(\cmd_mux_001|saved_grant[0]~q ),
	.always11(\router|always1~3_combout ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.mem_used_14(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest_generated(\sysid_qsys_0_control_slave_translator|av_waitrequest_generated~0_combout ),
	.wait_latency_counter_11(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~q ),
	.mem_used_15(mem_used_15),
	.Equal9(\router|Equal9~0_combout ),
	.av_waitrequest(av_waitrequest),
	.sink_ready1(\cmd_demux|sink_ready~7_combout ),
	.in_data_toggle(\crosser|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.Equal91(Equal9),
	.wait_latency_counter_12(\red_leds_s1_translator|wait_latency_counter[1]~1_combout ),
	.wait_latency_counter_0(\led_s1_translator|wait_latency_counter[0]~1_combout ),
	.WideOr0(\cmd_demux|WideOr0~7_combout ),
	.sink_ready2(sink_ready),
	.always12(\router|always1~5_combout ),
	.sink_ready3(\cmd_demux|sink_ready~12_combout ),
	.sink_ready4(\cmd_demux|sink_ready~13_combout ),
	.always13(\router|always1~6_combout ),
	.sink_ready5(\cmd_demux|sink_ready~14_combout ));

usb_system_usb_system_mm_interconnect_0_router_003_3 router_008(
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.always0(\router_008|always0~0_combout ));

endmodule

module usb_system_altera_avalon_sc_fifo (
	d_write,
	write_accepted,
	reset,
	read_latency_shift_reg_0,
	mem_67_0,
	mem_used_1,
	sink_ready,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
output 	mem_used_1;
input 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][67]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem[0][67]~1_combout ;
wire \mem_used[1]~0_combout ;


dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hB8FF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~1 (
	.dataa(\mem_used[0]~q ),
	.datab(sink_ready),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[0]~1_combout ),
	.cout());
defparam \mem_used[0]~1 .lut_mask = 16'hAFCF;
defparam \mem_used[0]~1 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_1),
	.datab(sink_ready),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hACFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_1 (
	reset,
	d_write,
	write_accepted,
	sink_in_reset,
	read_latency_shift_reg,
	out_valid,
	mem_67_0,
	full,
	mem_used_128,
	uav_read,
	m0_write,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	write_accepted;
input 	sink_in_reset;
input 	read_latency_shift_reg;
input 	out_valid;
output 	mem_67_0;
input 	full;
output 	mem_used_128;
input 	uav_read;
input 	m0_write;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[128][67]~q ;
wire \mem~254_combout ;
wire \write~0_combout ;
wire \mem_used~4_combout ;
wire \mem_used[127]~2_combout ;
wire \mem_used[127]~q ;
wire \mem_used~6_combout ;
wire \mem_used[126]~q ;
wire \mem_used~8_combout ;
wire \mem_used[125]~q ;
wire \mem_used~10_combout ;
wire \mem_used[124]~q ;
wire \mem_used~12_combout ;
wire \mem_used[123]~q ;
wire \mem_used~14_combout ;
wire \mem_used[122]~q ;
wire \mem_used~16_combout ;
wire \mem_used[121]~q ;
wire \mem_used~18_combout ;
wire \mem_used[120]~q ;
wire \mem_used~20_combout ;
wire \mem_used[119]~q ;
wire \mem_used~22_combout ;
wire \mem_used[118]~q ;
wire \mem_used~24_combout ;
wire \mem_used[117]~q ;
wire \mem_used~26_combout ;
wire \mem_used[116]~q ;
wire \mem_used~28_combout ;
wire \mem_used[115]~q ;
wire \mem_used~30_combout ;
wire \mem_used[114]~q ;
wire \mem_used~32_combout ;
wire \mem_used[113]~q ;
wire \mem_used~34_combout ;
wire \mem_used[112]~q ;
wire \mem_used~36_combout ;
wire \mem_used[111]~q ;
wire \mem_used~38_combout ;
wire \mem_used[110]~q ;
wire \mem_used~40_combout ;
wire \mem_used[109]~q ;
wire \mem_used~42_combout ;
wire \mem_used[108]~q ;
wire \mem_used~44_combout ;
wire \mem_used[107]~q ;
wire \mem_used~46_combout ;
wire \mem_used[106]~q ;
wire \mem_used~48_combout ;
wire \mem_used[105]~q ;
wire \mem_used~50_combout ;
wire \mem_used[104]~q ;
wire \mem_used~52_combout ;
wire \mem_used[103]~q ;
wire \mem_used~54_combout ;
wire \mem_used[102]~q ;
wire \mem_used~56_combout ;
wire \mem_used[101]~q ;
wire \mem_used~58_combout ;
wire \mem_used[100]~q ;
wire \mem_used~60_combout ;
wire \mem_used[99]~q ;
wire \mem_used~62_combout ;
wire \mem_used[98]~q ;
wire \mem_used~64_combout ;
wire \mem_used[97]~q ;
wire \mem_used~66_combout ;
wire \mem_used[96]~q ;
wire \mem_used~68_combout ;
wire \mem_used[95]~q ;
wire \mem_used~70_combout ;
wire \mem_used[94]~q ;
wire \mem_used~72_combout ;
wire \mem_used[93]~q ;
wire \mem_used~74_combout ;
wire \mem_used[92]~q ;
wire \mem_used~76_combout ;
wire \mem_used[91]~q ;
wire \mem_used~78_combout ;
wire \mem_used[90]~q ;
wire \mem_used~80_combout ;
wire \mem_used[89]~q ;
wire \mem_used~82_combout ;
wire \mem_used[88]~q ;
wire \mem_used~84_combout ;
wire \mem_used[87]~q ;
wire \mem_used~86_combout ;
wire \mem_used[86]~q ;
wire \mem_used~88_combout ;
wire \mem_used[85]~q ;
wire \mem_used~90_combout ;
wire \mem_used[84]~q ;
wire \mem_used~92_combout ;
wire \mem_used[83]~q ;
wire \mem_used~94_combout ;
wire \mem_used[82]~q ;
wire \mem_used~96_combout ;
wire \mem_used[81]~q ;
wire \mem_used~98_combout ;
wire \mem_used[80]~q ;
wire \mem_used~100_combout ;
wire \mem_used[79]~q ;
wire \mem_used~102_combout ;
wire \mem_used[78]~q ;
wire \mem_used~104_combout ;
wire \mem_used[77]~q ;
wire \mem_used~106_combout ;
wire \mem_used[76]~q ;
wire \mem_used~108_combout ;
wire \mem_used[75]~q ;
wire \mem_used~110_combout ;
wire \mem_used[74]~q ;
wire \mem_used~112_combout ;
wire \mem_used[73]~q ;
wire \mem_used~114_combout ;
wire \mem_used[72]~q ;
wire \mem_used~116_combout ;
wire \mem_used[71]~q ;
wire \mem_used~118_combout ;
wire \mem_used[70]~q ;
wire \mem_used~120_combout ;
wire \mem_used[69]~q ;
wire \mem_used~122_combout ;
wire \mem_used[68]~q ;
wire \mem_used~124_combout ;
wire \mem_used[67]~q ;
wire \mem_used~126_combout ;
wire \mem_used[66]~q ;
wire \mem_used~128_combout ;
wire \mem_used[65]~q ;
wire \mem_used~129_combout ;
wire \mem_used[64]~q ;
wire \mem_used~127_combout ;
wire \mem_used[63]~q ;
wire \mem_used~125_combout ;
wire \mem_used[62]~q ;
wire \mem_used~123_combout ;
wire \mem_used[61]~q ;
wire \mem_used~121_combout ;
wire \mem_used[60]~q ;
wire \mem_used~119_combout ;
wire \mem_used[59]~q ;
wire \mem_used~117_combout ;
wire \mem_used[58]~q ;
wire \mem_used~115_combout ;
wire \mem_used[57]~q ;
wire \mem_used~113_combout ;
wire \mem_used[56]~q ;
wire \mem_used~111_combout ;
wire \mem_used[55]~q ;
wire \mem_used~109_combout ;
wire \mem_used[54]~q ;
wire \mem_used~107_combout ;
wire \mem_used[53]~q ;
wire \mem_used~105_combout ;
wire \mem_used[52]~q ;
wire \mem_used~103_combout ;
wire \mem_used[51]~q ;
wire \mem_used~101_combout ;
wire \mem_used[50]~q ;
wire \mem_used~99_combout ;
wire \mem_used[49]~q ;
wire \mem_used~97_combout ;
wire \mem_used[48]~q ;
wire \mem_used~95_combout ;
wire \mem_used[47]~q ;
wire \mem_used~93_combout ;
wire \mem_used[46]~q ;
wire \mem_used~91_combout ;
wire \mem_used[45]~q ;
wire \mem_used~89_combout ;
wire \mem_used[44]~q ;
wire \mem_used~87_combout ;
wire \mem_used[43]~q ;
wire \mem_used~85_combout ;
wire \mem_used[42]~q ;
wire \mem_used~83_combout ;
wire \mem_used[41]~q ;
wire \mem_used~81_combout ;
wire \mem_used[40]~q ;
wire \mem_used~79_combout ;
wire \mem_used[39]~q ;
wire \mem_used~77_combout ;
wire \mem_used[38]~q ;
wire \mem_used~75_combout ;
wire \mem_used[37]~q ;
wire \mem_used~73_combout ;
wire \mem_used[36]~q ;
wire \mem_used~71_combout ;
wire \mem_used[35]~q ;
wire \mem_used~69_combout ;
wire \mem_used[34]~q ;
wire \mem_used~67_combout ;
wire \mem_used[33]~q ;
wire \mem_used~65_combout ;
wire \mem_used[32]~q ;
wire \mem_used~63_combout ;
wire \mem_used[31]~q ;
wire \mem_used~61_combout ;
wire \mem_used[30]~q ;
wire \mem_used~59_combout ;
wire \mem_used[29]~q ;
wire \mem_used~57_combout ;
wire \mem_used[28]~q ;
wire \mem_used~55_combout ;
wire \mem_used[27]~q ;
wire \mem_used~53_combout ;
wire \mem_used[26]~q ;
wire \mem_used~51_combout ;
wire \mem_used[25]~q ;
wire \mem_used~49_combout ;
wire \mem_used[24]~q ;
wire \mem_used~47_combout ;
wire \mem_used[23]~q ;
wire \mem_used~45_combout ;
wire \mem_used[22]~q ;
wire \mem_used~43_combout ;
wire \mem_used[21]~q ;
wire \mem_used~41_combout ;
wire \mem_used[20]~q ;
wire \mem_used~39_combout ;
wire \mem_used[19]~q ;
wire \mem_used~37_combout ;
wire \mem_used[18]~q ;
wire \mem_used~35_combout ;
wire \mem_used[17]~q ;
wire \mem_used~33_combout ;
wire \mem_used[16]~q ;
wire \mem_used~31_combout ;
wire \mem_used[15]~q ;
wire \mem_used~29_combout ;
wire \mem_used[14]~q ;
wire \mem_used~27_combout ;
wire \mem_used[13]~q ;
wire \mem_used~25_combout ;
wire \mem_used[12]~q ;
wire \mem_used~23_combout ;
wire \mem_used[11]~q ;
wire \mem_used~21_combout ;
wire \mem_used[10]~q ;
wire \mem_used~19_combout ;
wire \mem_used[9]~q ;
wire \mem_used~17_combout ;
wire \mem_used[8]~q ;
wire \mem_used~15_combout ;
wire \mem_used[7]~q ;
wire \mem_used~13_combout ;
wire \mem_used[6]~q ;
wire \mem_used~11_combout ;
wire \mem_used[5]~q ;
wire \mem_used~9_combout ;
wire \mem_used[4]~q ;
wire \mem_used~7_combout ;
wire \mem_used[3]~q ;
wire \mem_used~5_combout ;
wire \mem_used[2]~q ;
wire \mem_used~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \read~0_combout ;
wire \mem[127][67]~255_combout ;
wire \mem[127][67]~q ;
wire \mem[126][67]~252_combout ;
wire \mem[126][67]~253_combout ;
wire \mem[126][67]~q ;
wire \mem[125][67]~250_combout ;
wire \mem[125][67]~251_combout ;
wire \mem[125][67]~q ;
wire \mem[124][67]~248_combout ;
wire \mem[124][67]~249_combout ;
wire \mem[124][67]~q ;
wire \mem[123][67]~246_combout ;
wire \mem[123][67]~247_combout ;
wire \mem[123][67]~q ;
wire \mem[122][67]~244_combout ;
wire \mem[122][67]~245_combout ;
wire \mem[122][67]~q ;
wire \mem[121][67]~242_combout ;
wire \mem[121][67]~243_combout ;
wire \mem[121][67]~q ;
wire \mem[120][67]~240_combout ;
wire \mem[120][67]~241_combout ;
wire \mem[120][67]~q ;
wire \mem[119][67]~238_combout ;
wire \mem[119][67]~239_combout ;
wire \mem[119][67]~q ;
wire \mem[118][67]~236_combout ;
wire \mem[118][67]~237_combout ;
wire \mem[118][67]~q ;
wire \mem[117][67]~234_combout ;
wire \mem[117][67]~235_combout ;
wire \mem[117][67]~q ;
wire \mem[116][67]~232_combout ;
wire \mem[116][67]~233_combout ;
wire \mem[116][67]~q ;
wire \mem[115][67]~230_combout ;
wire \mem[115][67]~231_combout ;
wire \mem[115][67]~q ;
wire \mem[114][67]~228_combout ;
wire \mem[114][67]~229_combout ;
wire \mem[114][67]~q ;
wire \mem[113][67]~226_combout ;
wire \mem[113][67]~227_combout ;
wire \mem[113][67]~q ;
wire \mem[112][67]~224_combout ;
wire \mem[112][67]~225_combout ;
wire \mem[112][67]~q ;
wire \mem[111][67]~222_combout ;
wire \mem[111][67]~223_combout ;
wire \mem[111][67]~q ;
wire \mem[110][67]~220_combout ;
wire \mem[110][67]~221_combout ;
wire \mem[110][67]~q ;
wire \mem[109][67]~218_combout ;
wire \mem[109][67]~219_combout ;
wire \mem[109][67]~q ;
wire \mem[108][67]~216_combout ;
wire \mem[108][67]~217_combout ;
wire \mem[108][67]~q ;
wire \mem[107][67]~214_combout ;
wire \mem[107][67]~215_combout ;
wire \mem[107][67]~q ;
wire \mem[106][67]~212_combout ;
wire \mem[106][67]~213_combout ;
wire \mem[106][67]~q ;
wire \mem[105][67]~210_combout ;
wire \mem[105][67]~211_combout ;
wire \mem[105][67]~q ;
wire \mem[104][67]~208_combout ;
wire \mem[104][67]~209_combout ;
wire \mem[104][67]~q ;
wire \mem[103][67]~206_combout ;
wire \mem[103][67]~207_combout ;
wire \mem[103][67]~q ;
wire \mem[102][67]~204_combout ;
wire \mem[102][67]~205_combout ;
wire \mem[102][67]~q ;
wire \mem[101][67]~202_combout ;
wire \mem[101][67]~203_combout ;
wire \mem[101][67]~q ;
wire \mem[100][67]~200_combout ;
wire \mem[100][67]~201_combout ;
wire \mem[100][67]~q ;
wire \mem[99][67]~198_combout ;
wire \mem[99][67]~199_combout ;
wire \mem[99][67]~q ;
wire \mem[98][67]~196_combout ;
wire \mem[98][67]~197_combout ;
wire \mem[98][67]~q ;
wire \mem[97][67]~194_combout ;
wire \mem[97][67]~195_combout ;
wire \mem[97][67]~q ;
wire \mem[96][67]~192_combout ;
wire \mem[96][67]~193_combout ;
wire \mem[96][67]~q ;
wire \mem[95][67]~190_combout ;
wire \mem[95][67]~191_combout ;
wire \mem[95][67]~q ;
wire \mem[94][67]~188_combout ;
wire \mem[94][67]~189_combout ;
wire \mem[94][67]~q ;
wire \mem[93][67]~186_combout ;
wire \mem[93][67]~187_combout ;
wire \mem[93][67]~q ;
wire \mem[92][67]~184_combout ;
wire \mem[92][67]~185_combout ;
wire \mem[92][67]~q ;
wire \mem[91][67]~182_combout ;
wire \mem[91][67]~183_combout ;
wire \mem[91][67]~q ;
wire \mem[90][67]~180_combout ;
wire \mem[90][67]~181_combout ;
wire \mem[90][67]~q ;
wire \mem[89][67]~178_combout ;
wire \mem[89][67]~179_combout ;
wire \mem[89][67]~q ;
wire \mem[88][67]~176_combout ;
wire \mem[88][67]~177_combout ;
wire \mem[88][67]~q ;
wire \mem[87][67]~174_combout ;
wire \mem[87][67]~175_combout ;
wire \mem[87][67]~q ;
wire \mem[86][67]~172_combout ;
wire \mem[86][67]~173_combout ;
wire \mem[86][67]~q ;
wire \mem[85][67]~170_combout ;
wire \mem[85][67]~171_combout ;
wire \mem[85][67]~q ;
wire \mem[84][67]~168_combout ;
wire \mem[84][67]~169_combout ;
wire \mem[84][67]~q ;
wire \mem[83][67]~166_combout ;
wire \mem[83][67]~167_combout ;
wire \mem[83][67]~q ;
wire \mem[82][67]~164_combout ;
wire \mem[82][67]~165_combout ;
wire \mem[82][67]~q ;
wire \mem[81][67]~162_combout ;
wire \mem[81][67]~163_combout ;
wire \mem[81][67]~q ;
wire \mem[80][67]~160_combout ;
wire \mem[80][67]~161_combout ;
wire \mem[80][67]~q ;
wire \mem[79][67]~158_combout ;
wire \mem[79][67]~159_combout ;
wire \mem[79][67]~q ;
wire \mem[78][67]~156_combout ;
wire \mem[78][67]~157_combout ;
wire \mem[78][67]~q ;
wire \mem[77][67]~154_combout ;
wire \mem[77][67]~155_combout ;
wire \mem[77][67]~q ;
wire \mem[76][67]~152_combout ;
wire \mem[76][67]~153_combout ;
wire \mem[76][67]~q ;
wire \mem[75][67]~150_combout ;
wire \mem[75][67]~151_combout ;
wire \mem[75][67]~q ;
wire \mem[74][67]~148_combout ;
wire \mem[74][67]~149_combout ;
wire \mem[74][67]~q ;
wire \mem[73][67]~146_combout ;
wire \mem[73][67]~147_combout ;
wire \mem[73][67]~q ;
wire \mem[72][67]~144_combout ;
wire \mem[72][67]~145_combout ;
wire \mem[72][67]~q ;
wire \mem[71][67]~142_combout ;
wire \mem[71][67]~143_combout ;
wire \mem[71][67]~q ;
wire \mem[70][67]~140_combout ;
wire \mem[70][67]~141_combout ;
wire \mem[70][67]~q ;
wire \mem[69][67]~138_combout ;
wire \mem[69][67]~139_combout ;
wire \mem[69][67]~q ;
wire \mem[68][67]~136_combout ;
wire \mem[68][67]~137_combout ;
wire \mem[68][67]~q ;
wire \mem[67][67]~134_combout ;
wire \mem[67][67]~135_combout ;
wire \mem[67][67]~q ;
wire \mem[66][67]~132_combout ;
wire \mem[66][67]~133_combout ;
wire \mem[66][67]~q ;
wire \mem[65][67]~130_combout ;
wire \mem[65][67]~131_combout ;
wire \mem[65][67]~q ;
wire \mem[64][67]~128_combout ;
wire \mem[64][67]~129_combout ;
wire \mem[64][67]~q ;
wire \mem[63][67]~126_combout ;
wire \mem[63][67]~127_combout ;
wire \mem[63][67]~q ;
wire \mem[62][67]~124_combout ;
wire \mem[62][67]~125_combout ;
wire \mem[62][67]~q ;
wire \mem[61][67]~122_combout ;
wire \mem[61][67]~123_combout ;
wire \mem[61][67]~q ;
wire \mem[60][67]~120_combout ;
wire \mem[60][67]~121_combout ;
wire \mem[60][67]~q ;
wire \mem[59][67]~118_combout ;
wire \mem[59][67]~119_combout ;
wire \mem[59][67]~q ;
wire \mem[58][67]~116_combout ;
wire \mem[58][67]~117_combout ;
wire \mem[58][67]~q ;
wire \mem[57][67]~114_combout ;
wire \mem[57][67]~115_combout ;
wire \mem[57][67]~q ;
wire \mem[56][67]~112_combout ;
wire \mem[56][67]~113_combout ;
wire \mem[56][67]~q ;
wire \mem[55][67]~110_combout ;
wire \mem[55][67]~111_combout ;
wire \mem[55][67]~q ;
wire \mem[54][67]~108_combout ;
wire \mem[54][67]~109_combout ;
wire \mem[54][67]~q ;
wire \mem[53][67]~106_combout ;
wire \mem[53][67]~107_combout ;
wire \mem[53][67]~q ;
wire \mem[52][67]~104_combout ;
wire \mem[52][67]~105_combout ;
wire \mem[52][67]~q ;
wire \mem[51][67]~102_combout ;
wire \mem[51][67]~103_combout ;
wire \mem[51][67]~q ;
wire \mem[50][67]~100_combout ;
wire \mem[50][67]~101_combout ;
wire \mem[50][67]~q ;
wire \mem[49][67]~98_combout ;
wire \mem[49][67]~99_combout ;
wire \mem[49][67]~q ;
wire \mem[48][67]~96_combout ;
wire \mem[48][67]~97_combout ;
wire \mem[48][67]~q ;
wire \mem[47][67]~94_combout ;
wire \mem[47][67]~95_combout ;
wire \mem[47][67]~q ;
wire \mem[46][67]~92_combout ;
wire \mem[46][67]~93_combout ;
wire \mem[46][67]~q ;
wire \mem[45][67]~90_combout ;
wire \mem[45][67]~91_combout ;
wire \mem[45][67]~q ;
wire \mem[44][67]~88_combout ;
wire \mem[44][67]~89_combout ;
wire \mem[44][67]~q ;
wire \mem[43][67]~86_combout ;
wire \mem[43][67]~87_combout ;
wire \mem[43][67]~q ;
wire \mem[42][67]~84_combout ;
wire \mem[42][67]~85_combout ;
wire \mem[42][67]~q ;
wire \mem[41][67]~82_combout ;
wire \mem[41][67]~83_combout ;
wire \mem[41][67]~q ;
wire \mem[40][67]~80_combout ;
wire \mem[40][67]~81_combout ;
wire \mem[40][67]~q ;
wire \mem[39][67]~78_combout ;
wire \mem[39][67]~79_combout ;
wire \mem[39][67]~q ;
wire \mem[38][67]~76_combout ;
wire \mem[38][67]~77_combout ;
wire \mem[38][67]~q ;
wire \mem[37][67]~74_combout ;
wire \mem[37][67]~75_combout ;
wire \mem[37][67]~q ;
wire \mem[36][67]~72_combout ;
wire \mem[36][67]~73_combout ;
wire \mem[36][67]~q ;
wire \mem[35][67]~70_combout ;
wire \mem[35][67]~71_combout ;
wire \mem[35][67]~q ;
wire \mem[34][67]~68_combout ;
wire \mem[34][67]~69_combout ;
wire \mem[34][67]~q ;
wire \mem[33][67]~66_combout ;
wire \mem[33][67]~67_combout ;
wire \mem[33][67]~q ;
wire \mem[32][67]~64_combout ;
wire \mem[32][67]~65_combout ;
wire \mem[32][67]~q ;
wire \mem[31][67]~62_combout ;
wire \mem[31][67]~63_combout ;
wire \mem[31][67]~q ;
wire \mem[30][67]~60_combout ;
wire \mem[30][67]~61_combout ;
wire \mem[30][67]~q ;
wire \mem[29][67]~58_combout ;
wire \mem[29][67]~59_combout ;
wire \mem[29][67]~q ;
wire \mem[28][67]~56_combout ;
wire \mem[28][67]~57_combout ;
wire \mem[28][67]~q ;
wire \mem[27][67]~54_combout ;
wire \mem[27][67]~55_combout ;
wire \mem[27][67]~q ;
wire \mem[26][67]~52_combout ;
wire \mem[26][67]~53_combout ;
wire \mem[26][67]~q ;
wire \mem[25][67]~50_combout ;
wire \mem[25][67]~51_combout ;
wire \mem[25][67]~q ;
wire \mem[24][67]~48_combout ;
wire \mem[24][67]~49_combout ;
wire \mem[24][67]~q ;
wire \mem[23][67]~46_combout ;
wire \mem[23][67]~47_combout ;
wire \mem[23][67]~q ;
wire \mem[22][67]~44_combout ;
wire \mem[22][67]~45_combout ;
wire \mem[22][67]~q ;
wire \mem[21][67]~42_combout ;
wire \mem[21][67]~43_combout ;
wire \mem[21][67]~q ;
wire \mem[20][67]~40_combout ;
wire \mem[20][67]~41_combout ;
wire \mem[20][67]~q ;
wire \mem[19][67]~38_combout ;
wire \mem[19][67]~39_combout ;
wire \mem[19][67]~q ;
wire \mem[18][67]~36_combout ;
wire \mem[18][67]~37_combout ;
wire \mem[18][67]~q ;
wire \mem[17][67]~34_combout ;
wire \mem[17][67]~35_combout ;
wire \mem[17][67]~q ;
wire \mem[16][67]~32_combout ;
wire \mem[16][67]~33_combout ;
wire \mem[16][67]~q ;
wire \mem[15][67]~30_combout ;
wire \mem[15][67]~31_combout ;
wire \mem[15][67]~q ;
wire \mem[14][67]~28_combout ;
wire \mem[14][67]~29_combout ;
wire \mem[14][67]~q ;
wire \mem[13][67]~26_combout ;
wire \mem[13][67]~27_combout ;
wire \mem[13][67]~q ;
wire \mem[12][67]~24_combout ;
wire \mem[12][67]~25_combout ;
wire \mem[12][67]~q ;
wire \mem[11][67]~22_combout ;
wire \mem[11][67]~23_combout ;
wire \mem[11][67]~q ;
wire \mem[10][67]~20_combout ;
wire \mem[10][67]~21_combout ;
wire \mem[10][67]~q ;
wire \mem[9][67]~18_combout ;
wire \mem[9][67]~19_combout ;
wire \mem[9][67]~q ;
wire \mem[8][67]~16_combout ;
wire \mem[8][67]~17_combout ;
wire \mem[8][67]~q ;
wire \mem[7][67]~14_combout ;
wire \mem[7][67]~15_combout ;
wire \mem[7][67]~q ;
wire \mem[6][67]~12_combout ;
wire \mem[6][67]~13_combout ;
wire \mem[6][67]~q ;
wire \mem[5][67]~10_combout ;
wire \mem[5][67]~11_combout ;
wire \mem[5][67]~q ;
wire \mem[4][67]~8_combout ;
wire \mem[4][67]~9_combout ;
wire \mem[4][67]~q ;
wire \mem[3][67]~6_combout ;
wire \mem[3][67]~7_combout ;
wire \mem[3][67]~q ;
wire \mem[2][67]~4_combout ;
wire \mem[2][67]~5_combout ;
wire \mem[2][67]~q ;
wire \mem[1][67]~2_combout ;
wire \mem[1][67]~3_combout ;
wire \mem[1][67]~q ;
wire \mem[0][67]~0_combout ;
wire \mem[0][67]~1_combout ;
wire \mem_used[128]~0_combout ;


dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[128] (
	.clk(clk),
	.d(\mem_used[128]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_128),
	.prn(vcc));
defparam \mem_used[128] .is_wysiwyg = "true";
defparam \mem_used[128] .power_up = "low";

dffeas \mem[128][67] (
	.clk(clk),
	.d(\mem~254_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[128][67]~q ),
	.prn(vcc));
defparam \mem[128][67] .is_wysiwyg = "true";
defparam \mem[128][67] .power_up = "low";

cycloneive_lcell_comb \mem~254 (
	.dataa(\mem[128][67]~q ),
	.datab(mem_used_128),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~254_combout ),
	.cout());
defparam \mem~254 .lut_mask = 16'hB8FF;
defparam \mem~254 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~0 (
	.dataa(sink_in_reset),
	.datab(uav_read),
	.datac(m0_write),
	.datad(full),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFEFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used~4 (
	.dataa(mem_used_128),
	.datab(\write~0_combout ),
	.datac(\mem_used[126]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used~4_combout ),
	.cout());
defparam \mem_used~4 .lut_mask = 16'hFEFE;
defparam \mem_used~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[127]~2 (
	.dataa(\read~0_combout ),
	.datab(full),
	.datac(read_latency_shift_reg),
	.datad(m0_write),
	.cin(gnd),
	.combout(\mem_used[127]~2_combout ),
	.cout());
defparam \mem_used[127]~2 .lut_mask = 16'h6996;
defparam \mem_used[127]~2 .sum_lutc_input = "datac";

dffeas \mem_used[127] (
	.clk(clk),
	.d(\mem_used~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[127]~q ),
	.prn(vcc));
defparam \mem_used[127] .is_wysiwyg = "true";
defparam \mem_used[127] .power_up = "low";

cycloneive_lcell_comb \mem_used~6 (
	.dataa(\mem_used[125]~q ),
	.datab(\mem_used[127]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~6_combout ),
	.cout());
defparam \mem_used~6 .lut_mask = 16'hAACC;
defparam \mem_used~6 .sum_lutc_input = "datac";

dffeas \mem_used[126] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[126]~q ),
	.prn(vcc));
defparam \mem_used[126] .is_wysiwyg = "true";
defparam \mem_used[126] .power_up = "low";

cycloneive_lcell_comb \mem_used~8 (
	.dataa(\mem_used[124]~q ),
	.datab(\mem_used[126]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~8_combout ),
	.cout());
defparam \mem_used~8 .lut_mask = 16'hAACC;
defparam \mem_used~8 .sum_lutc_input = "datac";

dffeas \mem_used[125] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[125]~q ),
	.prn(vcc));
defparam \mem_used[125] .is_wysiwyg = "true";
defparam \mem_used[125] .power_up = "low";

cycloneive_lcell_comb \mem_used~10 (
	.dataa(\mem_used[123]~q ),
	.datab(\mem_used[125]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~10_combout ),
	.cout());
defparam \mem_used~10 .lut_mask = 16'hAACC;
defparam \mem_used~10 .sum_lutc_input = "datac";

dffeas \mem_used[124] (
	.clk(clk),
	.d(\mem_used~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[124]~q ),
	.prn(vcc));
defparam \mem_used[124] .is_wysiwyg = "true";
defparam \mem_used[124] .power_up = "low";

cycloneive_lcell_comb \mem_used~12 (
	.dataa(\mem_used[122]~q ),
	.datab(\mem_used[124]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~12_combout ),
	.cout());
defparam \mem_used~12 .lut_mask = 16'hAACC;
defparam \mem_used~12 .sum_lutc_input = "datac";

dffeas \mem_used[123] (
	.clk(clk),
	.d(\mem_used~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[123]~q ),
	.prn(vcc));
defparam \mem_used[123] .is_wysiwyg = "true";
defparam \mem_used[123] .power_up = "low";

cycloneive_lcell_comb \mem_used~14 (
	.dataa(\mem_used[121]~q ),
	.datab(\mem_used[123]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~14_combout ),
	.cout());
defparam \mem_used~14 .lut_mask = 16'hAACC;
defparam \mem_used~14 .sum_lutc_input = "datac";

dffeas \mem_used[122] (
	.clk(clk),
	.d(\mem_used~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[122]~q ),
	.prn(vcc));
defparam \mem_used[122] .is_wysiwyg = "true";
defparam \mem_used[122] .power_up = "low";

cycloneive_lcell_comb \mem_used~16 (
	.dataa(\mem_used[120]~q ),
	.datab(\mem_used[122]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~16_combout ),
	.cout());
defparam \mem_used~16 .lut_mask = 16'hAACC;
defparam \mem_used~16 .sum_lutc_input = "datac";

dffeas \mem_used[121] (
	.clk(clk),
	.d(\mem_used~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[121]~q ),
	.prn(vcc));
defparam \mem_used[121] .is_wysiwyg = "true";
defparam \mem_used[121] .power_up = "low";

cycloneive_lcell_comb \mem_used~18 (
	.dataa(\mem_used[119]~q ),
	.datab(\mem_used[121]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~18_combout ),
	.cout());
defparam \mem_used~18 .lut_mask = 16'hAACC;
defparam \mem_used~18 .sum_lutc_input = "datac";

dffeas \mem_used[120] (
	.clk(clk),
	.d(\mem_used~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[120]~q ),
	.prn(vcc));
defparam \mem_used[120] .is_wysiwyg = "true";
defparam \mem_used[120] .power_up = "low";

cycloneive_lcell_comb \mem_used~20 (
	.dataa(\mem_used[118]~q ),
	.datab(\mem_used[120]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~20_combout ),
	.cout());
defparam \mem_used~20 .lut_mask = 16'hAACC;
defparam \mem_used~20 .sum_lutc_input = "datac";

dffeas \mem_used[119] (
	.clk(clk),
	.d(\mem_used~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[119]~q ),
	.prn(vcc));
defparam \mem_used[119] .is_wysiwyg = "true";
defparam \mem_used[119] .power_up = "low";

cycloneive_lcell_comb \mem_used~22 (
	.dataa(\mem_used[117]~q ),
	.datab(\mem_used[119]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~22_combout ),
	.cout());
defparam \mem_used~22 .lut_mask = 16'hAACC;
defparam \mem_used~22 .sum_lutc_input = "datac";

dffeas \mem_used[118] (
	.clk(clk),
	.d(\mem_used~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[118]~q ),
	.prn(vcc));
defparam \mem_used[118] .is_wysiwyg = "true";
defparam \mem_used[118] .power_up = "low";

cycloneive_lcell_comb \mem_used~24 (
	.dataa(\mem_used[116]~q ),
	.datab(\mem_used[118]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~24_combout ),
	.cout());
defparam \mem_used~24 .lut_mask = 16'hAACC;
defparam \mem_used~24 .sum_lutc_input = "datac";

dffeas \mem_used[117] (
	.clk(clk),
	.d(\mem_used~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[117]~q ),
	.prn(vcc));
defparam \mem_used[117] .is_wysiwyg = "true";
defparam \mem_used[117] .power_up = "low";

cycloneive_lcell_comb \mem_used~26 (
	.dataa(\mem_used[115]~q ),
	.datab(\mem_used[117]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~26_combout ),
	.cout());
defparam \mem_used~26 .lut_mask = 16'hAACC;
defparam \mem_used~26 .sum_lutc_input = "datac";

dffeas \mem_used[116] (
	.clk(clk),
	.d(\mem_used~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[116]~q ),
	.prn(vcc));
defparam \mem_used[116] .is_wysiwyg = "true";
defparam \mem_used[116] .power_up = "low";

cycloneive_lcell_comb \mem_used~28 (
	.dataa(\mem_used[114]~q ),
	.datab(\mem_used[116]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~28_combout ),
	.cout());
defparam \mem_used~28 .lut_mask = 16'hAACC;
defparam \mem_used~28 .sum_lutc_input = "datac";

dffeas \mem_used[115] (
	.clk(clk),
	.d(\mem_used~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[115]~q ),
	.prn(vcc));
defparam \mem_used[115] .is_wysiwyg = "true";
defparam \mem_used[115] .power_up = "low";

cycloneive_lcell_comb \mem_used~30 (
	.dataa(\mem_used[113]~q ),
	.datab(\mem_used[115]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~30_combout ),
	.cout());
defparam \mem_used~30 .lut_mask = 16'hAACC;
defparam \mem_used~30 .sum_lutc_input = "datac";

dffeas \mem_used[114] (
	.clk(clk),
	.d(\mem_used~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[114]~q ),
	.prn(vcc));
defparam \mem_used[114] .is_wysiwyg = "true";
defparam \mem_used[114] .power_up = "low";

cycloneive_lcell_comb \mem_used~32 (
	.dataa(\mem_used[112]~q ),
	.datab(\mem_used[114]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~32_combout ),
	.cout());
defparam \mem_used~32 .lut_mask = 16'hAACC;
defparam \mem_used~32 .sum_lutc_input = "datac";

dffeas \mem_used[113] (
	.clk(clk),
	.d(\mem_used~32_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[113]~q ),
	.prn(vcc));
defparam \mem_used[113] .is_wysiwyg = "true";
defparam \mem_used[113] .power_up = "low";

cycloneive_lcell_comb \mem_used~34 (
	.dataa(\mem_used[111]~q ),
	.datab(\mem_used[113]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~34_combout ),
	.cout());
defparam \mem_used~34 .lut_mask = 16'hAACC;
defparam \mem_used~34 .sum_lutc_input = "datac";

dffeas \mem_used[112] (
	.clk(clk),
	.d(\mem_used~34_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[112]~q ),
	.prn(vcc));
defparam \mem_used[112] .is_wysiwyg = "true";
defparam \mem_used[112] .power_up = "low";

cycloneive_lcell_comb \mem_used~36 (
	.dataa(\mem_used[110]~q ),
	.datab(\mem_used[112]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~36_combout ),
	.cout());
defparam \mem_used~36 .lut_mask = 16'hAACC;
defparam \mem_used~36 .sum_lutc_input = "datac";

dffeas \mem_used[111] (
	.clk(clk),
	.d(\mem_used~36_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[111]~q ),
	.prn(vcc));
defparam \mem_used[111] .is_wysiwyg = "true";
defparam \mem_used[111] .power_up = "low";

cycloneive_lcell_comb \mem_used~38 (
	.dataa(\mem_used[109]~q ),
	.datab(\mem_used[111]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~38_combout ),
	.cout());
defparam \mem_used~38 .lut_mask = 16'hAACC;
defparam \mem_used~38 .sum_lutc_input = "datac";

dffeas \mem_used[110] (
	.clk(clk),
	.d(\mem_used~38_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[110]~q ),
	.prn(vcc));
defparam \mem_used[110] .is_wysiwyg = "true";
defparam \mem_used[110] .power_up = "low";

cycloneive_lcell_comb \mem_used~40 (
	.dataa(\mem_used[108]~q ),
	.datab(\mem_used[110]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~40_combout ),
	.cout());
defparam \mem_used~40 .lut_mask = 16'hAACC;
defparam \mem_used~40 .sum_lutc_input = "datac";

dffeas \mem_used[109] (
	.clk(clk),
	.d(\mem_used~40_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[109]~q ),
	.prn(vcc));
defparam \mem_used[109] .is_wysiwyg = "true";
defparam \mem_used[109] .power_up = "low";

cycloneive_lcell_comb \mem_used~42 (
	.dataa(\mem_used[107]~q ),
	.datab(\mem_used[109]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~42_combout ),
	.cout());
defparam \mem_used~42 .lut_mask = 16'hAACC;
defparam \mem_used~42 .sum_lutc_input = "datac";

dffeas \mem_used[108] (
	.clk(clk),
	.d(\mem_used~42_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[108]~q ),
	.prn(vcc));
defparam \mem_used[108] .is_wysiwyg = "true";
defparam \mem_used[108] .power_up = "low";

cycloneive_lcell_comb \mem_used~44 (
	.dataa(\mem_used[106]~q ),
	.datab(\mem_used[108]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~44_combout ),
	.cout());
defparam \mem_used~44 .lut_mask = 16'hAACC;
defparam \mem_used~44 .sum_lutc_input = "datac";

dffeas \mem_used[107] (
	.clk(clk),
	.d(\mem_used~44_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[107]~q ),
	.prn(vcc));
defparam \mem_used[107] .is_wysiwyg = "true";
defparam \mem_used[107] .power_up = "low";

cycloneive_lcell_comb \mem_used~46 (
	.dataa(\mem_used[105]~q ),
	.datab(\mem_used[107]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~46_combout ),
	.cout());
defparam \mem_used~46 .lut_mask = 16'hAACC;
defparam \mem_used~46 .sum_lutc_input = "datac";

dffeas \mem_used[106] (
	.clk(clk),
	.d(\mem_used~46_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[106]~q ),
	.prn(vcc));
defparam \mem_used[106] .is_wysiwyg = "true";
defparam \mem_used[106] .power_up = "low";

cycloneive_lcell_comb \mem_used~48 (
	.dataa(\mem_used[104]~q ),
	.datab(\mem_used[106]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~48_combout ),
	.cout());
defparam \mem_used~48 .lut_mask = 16'hAACC;
defparam \mem_used~48 .sum_lutc_input = "datac";

dffeas \mem_used[105] (
	.clk(clk),
	.d(\mem_used~48_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[105]~q ),
	.prn(vcc));
defparam \mem_used[105] .is_wysiwyg = "true";
defparam \mem_used[105] .power_up = "low";

cycloneive_lcell_comb \mem_used~50 (
	.dataa(\mem_used[103]~q ),
	.datab(\mem_used[105]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~50_combout ),
	.cout());
defparam \mem_used~50 .lut_mask = 16'hAACC;
defparam \mem_used~50 .sum_lutc_input = "datac";

dffeas \mem_used[104] (
	.clk(clk),
	.d(\mem_used~50_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[104]~q ),
	.prn(vcc));
defparam \mem_used[104] .is_wysiwyg = "true";
defparam \mem_used[104] .power_up = "low";

cycloneive_lcell_comb \mem_used~52 (
	.dataa(\mem_used[102]~q ),
	.datab(\mem_used[104]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~52_combout ),
	.cout());
defparam \mem_used~52 .lut_mask = 16'hAACC;
defparam \mem_used~52 .sum_lutc_input = "datac";

dffeas \mem_used[103] (
	.clk(clk),
	.d(\mem_used~52_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[103]~q ),
	.prn(vcc));
defparam \mem_used[103] .is_wysiwyg = "true";
defparam \mem_used[103] .power_up = "low";

cycloneive_lcell_comb \mem_used~54 (
	.dataa(\mem_used[101]~q ),
	.datab(\mem_used[103]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~54_combout ),
	.cout());
defparam \mem_used~54 .lut_mask = 16'hAACC;
defparam \mem_used~54 .sum_lutc_input = "datac";

dffeas \mem_used[102] (
	.clk(clk),
	.d(\mem_used~54_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[102]~q ),
	.prn(vcc));
defparam \mem_used[102] .is_wysiwyg = "true";
defparam \mem_used[102] .power_up = "low";

cycloneive_lcell_comb \mem_used~56 (
	.dataa(\mem_used[100]~q ),
	.datab(\mem_used[102]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~56_combout ),
	.cout());
defparam \mem_used~56 .lut_mask = 16'hAACC;
defparam \mem_used~56 .sum_lutc_input = "datac";

dffeas \mem_used[101] (
	.clk(clk),
	.d(\mem_used~56_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[101]~q ),
	.prn(vcc));
defparam \mem_used[101] .is_wysiwyg = "true";
defparam \mem_used[101] .power_up = "low";

cycloneive_lcell_comb \mem_used~58 (
	.dataa(\mem_used[99]~q ),
	.datab(\mem_used[101]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~58_combout ),
	.cout());
defparam \mem_used~58 .lut_mask = 16'hAACC;
defparam \mem_used~58 .sum_lutc_input = "datac";

dffeas \mem_used[100] (
	.clk(clk),
	.d(\mem_used~58_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[100]~q ),
	.prn(vcc));
defparam \mem_used[100] .is_wysiwyg = "true";
defparam \mem_used[100] .power_up = "low";

cycloneive_lcell_comb \mem_used~60 (
	.dataa(\mem_used[98]~q ),
	.datab(\mem_used[100]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~60_combout ),
	.cout());
defparam \mem_used~60 .lut_mask = 16'hAACC;
defparam \mem_used~60 .sum_lutc_input = "datac";

dffeas \mem_used[99] (
	.clk(clk),
	.d(\mem_used~60_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[99]~q ),
	.prn(vcc));
defparam \mem_used[99] .is_wysiwyg = "true";
defparam \mem_used[99] .power_up = "low";

cycloneive_lcell_comb \mem_used~62 (
	.dataa(\mem_used[97]~q ),
	.datab(\mem_used[99]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~62_combout ),
	.cout());
defparam \mem_used~62 .lut_mask = 16'hAACC;
defparam \mem_used~62 .sum_lutc_input = "datac";

dffeas \mem_used[98] (
	.clk(clk),
	.d(\mem_used~62_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[98]~q ),
	.prn(vcc));
defparam \mem_used[98] .is_wysiwyg = "true";
defparam \mem_used[98] .power_up = "low";

cycloneive_lcell_comb \mem_used~64 (
	.dataa(\mem_used[96]~q ),
	.datab(\mem_used[98]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~64_combout ),
	.cout());
defparam \mem_used~64 .lut_mask = 16'hAACC;
defparam \mem_used~64 .sum_lutc_input = "datac";

dffeas \mem_used[97] (
	.clk(clk),
	.d(\mem_used~64_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[97]~q ),
	.prn(vcc));
defparam \mem_used[97] .is_wysiwyg = "true";
defparam \mem_used[97] .power_up = "low";

cycloneive_lcell_comb \mem_used~66 (
	.dataa(\mem_used[95]~q ),
	.datab(\mem_used[97]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~66_combout ),
	.cout());
defparam \mem_used~66 .lut_mask = 16'hAACC;
defparam \mem_used~66 .sum_lutc_input = "datac";

dffeas \mem_used[96] (
	.clk(clk),
	.d(\mem_used~66_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[96]~q ),
	.prn(vcc));
defparam \mem_used[96] .is_wysiwyg = "true";
defparam \mem_used[96] .power_up = "low";

cycloneive_lcell_comb \mem_used~68 (
	.dataa(\mem_used[94]~q ),
	.datab(\mem_used[96]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~68_combout ),
	.cout());
defparam \mem_used~68 .lut_mask = 16'hAACC;
defparam \mem_used~68 .sum_lutc_input = "datac";

dffeas \mem_used[95] (
	.clk(clk),
	.d(\mem_used~68_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[95]~q ),
	.prn(vcc));
defparam \mem_used[95] .is_wysiwyg = "true";
defparam \mem_used[95] .power_up = "low";

cycloneive_lcell_comb \mem_used~70 (
	.dataa(\mem_used[93]~q ),
	.datab(\mem_used[95]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~70_combout ),
	.cout());
defparam \mem_used~70 .lut_mask = 16'hAACC;
defparam \mem_used~70 .sum_lutc_input = "datac";

dffeas \mem_used[94] (
	.clk(clk),
	.d(\mem_used~70_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[94]~q ),
	.prn(vcc));
defparam \mem_used[94] .is_wysiwyg = "true";
defparam \mem_used[94] .power_up = "low";

cycloneive_lcell_comb \mem_used~72 (
	.dataa(\mem_used[92]~q ),
	.datab(\mem_used[94]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~72_combout ),
	.cout());
defparam \mem_used~72 .lut_mask = 16'hAACC;
defparam \mem_used~72 .sum_lutc_input = "datac";

dffeas \mem_used[93] (
	.clk(clk),
	.d(\mem_used~72_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[93]~q ),
	.prn(vcc));
defparam \mem_used[93] .is_wysiwyg = "true";
defparam \mem_used[93] .power_up = "low";

cycloneive_lcell_comb \mem_used~74 (
	.dataa(\mem_used[91]~q ),
	.datab(\mem_used[93]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~74_combout ),
	.cout());
defparam \mem_used~74 .lut_mask = 16'hAACC;
defparam \mem_used~74 .sum_lutc_input = "datac";

dffeas \mem_used[92] (
	.clk(clk),
	.d(\mem_used~74_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[92]~q ),
	.prn(vcc));
defparam \mem_used[92] .is_wysiwyg = "true";
defparam \mem_used[92] .power_up = "low";

cycloneive_lcell_comb \mem_used~76 (
	.dataa(\mem_used[90]~q ),
	.datab(\mem_used[92]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~76_combout ),
	.cout());
defparam \mem_used~76 .lut_mask = 16'hAACC;
defparam \mem_used~76 .sum_lutc_input = "datac";

dffeas \mem_used[91] (
	.clk(clk),
	.d(\mem_used~76_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[91]~q ),
	.prn(vcc));
defparam \mem_used[91] .is_wysiwyg = "true";
defparam \mem_used[91] .power_up = "low";

cycloneive_lcell_comb \mem_used~78 (
	.dataa(\mem_used[89]~q ),
	.datab(\mem_used[91]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~78_combout ),
	.cout());
defparam \mem_used~78 .lut_mask = 16'hAACC;
defparam \mem_used~78 .sum_lutc_input = "datac";

dffeas \mem_used[90] (
	.clk(clk),
	.d(\mem_used~78_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[90]~q ),
	.prn(vcc));
defparam \mem_used[90] .is_wysiwyg = "true";
defparam \mem_used[90] .power_up = "low";

cycloneive_lcell_comb \mem_used~80 (
	.dataa(\mem_used[88]~q ),
	.datab(\mem_used[90]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~80_combout ),
	.cout());
defparam \mem_used~80 .lut_mask = 16'hAACC;
defparam \mem_used~80 .sum_lutc_input = "datac";

dffeas \mem_used[89] (
	.clk(clk),
	.d(\mem_used~80_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[89]~q ),
	.prn(vcc));
defparam \mem_used[89] .is_wysiwyg = "true";
defparam \mem_used[89] .power_up = "low";

cycloneive_lcell_comb \mem_used~82 (
	.dataa(\mem_used[87]~q ),
	.datab(\mem_used[89]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~82_combout ),
	.cout());
defparam \mem_used~82 .lut_mask = 16'hAACC;
defparam \mem_used~82 .sum_lutc_input = "datac";

dffeas \mem_used[88] (
	.clk(clk),
	.d(\mem_used~82_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[88]~q ),
	.prn(vcc));
defparam \mem_used[88] .is_wysiwyg = "true";
defparam \mem_used[88] .power_up = "low";

cycloneive_lcell_comb \mem_used~84 (
	.dataa(\mem_used[86]~q ),
	.datab(\mem_used[88]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~84_combout ),
	.cout());
defparam \mem_used~84 .lut_mask = 16'hAACC;
defparam \mem_used~84 .sum_lutc_input = "datac";

dffeas \mem_used[87] (
	.clk(clk),
	.d(\mem_used~84_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[87]~q ),
	.prn(vcc));
defparam \mem_used[87] .is_wysiwyg = "true";
defparam \mem_used[87] .power_up = "low";

cycloneive_lcell_comb \mem_used~86 (
	.dataa(\mem_used[85]~q ),
	.datab(\mem_used[87]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~86_combout ),
	.cout());
defparam \mem_used~86 .lut_mask = 16'hAACC;
defparam \mem_used~86 .sum_lutc_input = "datac";

dffeas \mem_used[86] (
	.clk(clk),
	.d(\mem_used~86_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[86]~q ),
	.prn(vcc));
defparam \mem_used[86] .is_wysiwyg = "true";
defparam \mem_used[86] .power_up = "low";

cycloneive_lcell_comb \mem_used~88 (
	.dataa(\mem_used[84]~q ),
	.datab(\mem_used[86]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~88_combout ),
	.cout());
defparam \mem_used~88 .lut_mask = 16'hAACC;
defparam \mem_used~88 .sum_lutc_input = "datac";

dffeas \mem_used[85] (
	.clk(clk),
	.d(\mem_used~88_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[85]~q ),
	.prn(vcc));
defparam \mem_used[85] .is_wysiwyg = "true";
defparam \mem_used[85] .power_up = "low";

cycloneive_lcell_comb \mem_used~90 (
	.dataa(\mem_used[83]~q ),
	.datab(\mem_used[85]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~90_combout ),
	.cout());
defparam \mem_used~90 .lut_mask = 16'hAACC;
defparam \mem_used~90 .sum_lutc_input = "datac";

dffeas \mem_used[84] (
	.clk(clk),
	.d(\mem_used~90_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[84]~q ),
	.prn(vcc));
defparam \mem_used[84] .is_wysiwyg = "true";
defparam \mem_used[84] .power_up = "low";

cycloneive_lcell_comb \mem_used~92 (
	.dataa(\mem_used[82]~q ),
	.datab(\mem_used[84]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~92_combout ),
	.cout());
defparam \mem_used~92 .lut_mask = 16'hAACC;
defparam \mem_used~92 .sum_lutc_input = "datac";

dffeas \mem_used[83] (
	.clk(clk),
	.d(\mem_used~92_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[83]~q ),
	.prn(vcc));
defparam \mem_used[83] .is_wysiwyg = "true";
defparam \mem_used[83] .power_up = "low";

cycloneive_lcell_comb \mem_used~94 (
	.dataa(\mem_used[81]~q ),
	.datab(\mem_used[83]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~94_combout ),
	.cout());
defparam \mem_used~94 .lut_mask = 16'hAACC;
defparam \mem_used~94 .sum_lutc_input = "datac";

dffeas \mem_used[82] (
	.clk(clk),
	.d(\mem_used~94_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[82]~q ),
	.prn(vcc));
defparam \mem_used[82] .is_wysiwyg = "true";
defparam \mem_used[82] .power_up = "low";

cycloneive_lcell_comb \mem_used~96 (
	.dataa(\mem_used[80]~q ),
	.datab(\mem_used[82]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~96_combout ),
	.cout());
defparam \mem_used~96 .lut_mask = 16'hAACC;
defparam \mem_used~96 .sum_lutc_input = "datac";

dffeas \mem_used[81] (
	.clk(clk),
	.d(\mem_used~96_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[81]~q ),
	.prn(vcc));
defparam \mem_used[81] .is_wysiwyg = "true";
defparam \mem_used[81] .power_up = "low";

cycloneive_lcell_comb \mem_used~98 (
	.dataa(\mem_used[79]~q ),
	.datab(\mem_used[81]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~98_combout ),
	.cout());
defparam \mem_used~98 .lut_mask = 16'hAACC;
defparam \mem_used~98 .sum_lutc_input = "datac";

dffeas \mem_used[80] (
	.clk(clk),
	.d(\mem_used~98_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[80]~q ),
	.prn(vcc));
defparam \mem_used[80] .is_wysiwyg = "true";
defparam \mem_used[80] .power_up = "low";

cycloneive_lcell_comb \mem_used~100 (
	.dataa(\mem_used[78]~q ),
	.datab(\mem_used[80]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~100_combout ),
	.cout());
defparam \mem_used~100 .lut_mask = 16'hAACC;
defparam \mem_used~100 .sum_lutc_input = "datac";

dffeas \mem_used[79] (
	.clk(clk),
	.d(\mem_used~100_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[79]~q ),
	.prn(vcc));
defparam \mem_used[79] .is_wysiwyg = "true";
defparam \mem_used[79] .power_up = "low";

cycloneive_lcell_comb \mem_used~102 (
	.dataa(\mem_used[77]~q ),
	.datab(\mem_used[79]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~102_combout ),
	.cout());
defparam \mem_used~102 .lut_mask = 16'hAACC;
defparam \mem_used~102 .sum_lutc_input = "datac";

dffeas \mem_used[78] (
	.clk(clk),
	.d(\mem_used~102_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[78]~q ),
	.prn(vcc));
defparam \mem_used[78] .is_wysiwyg = "true";
defparam \mem_used[78] .power_up = "low";

cycloneive_lcell_comb \mem_used~104 (
	.dataa(\mem_used[76]~q ),
	.datab(\mem_used[78]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~104_combout ),
	.cout());
defparam \mem_used~104 .lut_mask = 16'hAACC;
defparam \mem_used~104 .sum_lutc_input = "datac";

dffeas \mem_used[77] (
	.clk(clk),
	.d(\mem_used~104_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[77]~q ),
	.prn(vcc));
defparam \mem_used[77] .is_wysiwyg = "true";
defparam \mem_used[77] .power_up = "low";

cycloneive_lcell_comb \mem_used~106 (
	.dataa(\mem_used[75]~q ),
	.datab(\mem_used[77]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~106_combout ),
	.cout());
defparam \mem_used~106 .lut_mask = 16'hAACC;
defparam \mem_used~106 .sum_lutc_input = "datac";

dffeas \mem_used[76] (
	.clk(clk),
	.d(\mem_used~106_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[76]~q ),
	.prn(vcc));
defparam \mem_used[76] .is_wysiwyg = "true";
defparam \mem_used[76] .power_up = "low";

cycloneive_lcell_comb \mem_used~108 (
	.dataa(\mem_used[74]~q ),
	.datab(\mem_used[76]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~108_combout ),
	.cout());
defparam \mem_used~108 .lut_mask = 16'hAACC;
defparam \mem_used~108 .sum_lutc_input = "datac";

dffeas \mem_used[75] (
	.clk(clk),
	.d(\mem_used~108_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[75]~q ),
	.prn(vcc));
defparam \mem_used[75] .is_wysiwyg = "true";
defparam \mem_used[75] .power_up = "low";

cycloneive_lcell_comb \mem_used~110 (
	.dataa(\mem_used[73]~q ),
	.datab(\mem_used[75]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~110_combout ),
	.cout());
defparam \mem_used~110 .lut_mask = 16'hAACC;
defparam \mem_used~110 .sum_lutc_input = "datac";

dffeas \mem_used[74] (
	.clk(clk),
	.d(\mem_used~110_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[74]~q ),
	.prn(vcc));
defparam \mem_used[74] .is_wysiwyg = "true";
defparam \mem_used[74] .power_up = "low";

cycloneive_lcell_comb \mem_used~112 (
	.dataa(\mem_used[72]~q ),
	.datab(\mem_used[74]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~112_combout ),
	.cout());
defparam \mem_used~112 .lut_mask = 16'hAACC;
defparam \mem_used~112 .sum_lutc_input = "datac";

dffeas \mem_used[73] (
	.clk(clk),
	.d(\mem_used~112_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[73]~q ),
	.prn(vcc));
defparam \mem_used[73] .is_wysiwyg = "true";
defparam \mem_used[73] .power_up = "low";

cycloneive_lcell_comb \mem_used~114 (
	.dataa(\mem_used[71]~q ),
	.datab(\mem_used[73]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~114_combout ),
	.cout());
defparam \mem_used~114 .lut_mask = 16'hAACC;
defparam \mem_used~114 .sum_lutc_input = "datac";

dffeas \mem_used[72] (
	.clk(clk),
	.d(\mem_used~114_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[72]~q ),
	.prn(vcc));
defparam \mem_used[72] .is_wysiwyg = "true";
defparam \mem_used[72] .power_up = "low";

cycloneive_lcell_comb \mem_used~116 (
	.dataa(\mem_used[70]~q ),
	.datab(\mem_used[72]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~116_combout ),
	.cout());
defparam \mem_used~116 .lut_mask = 16'hAACC;
defparam \mem_used~116 .sum_lutc_input = "datac";

dffeas \mem_used[71] (
	.clk(clk),
	.d(\mem_used~116_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[71]~q ),
	.prn(vcc));
defparam \mem_used[71] .is_wysiwyg = "true";
defparam \mem_used[71] .power_up = "low";

cycloneive_lcell_comb \mem_used~118 (
	.dataa(\mem_used[69]~q ),
	.datab(\mem_used[71]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~118_combout ),
	.cout());
defparam \mem_used~118 .lut_mask = 16'hAACC;
defparam \mem_used~118 .sum_lutc_input = "datac";

dffeas \mem_used[70] (
	.clk(clk),
	.d(\mem_used~118_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[70]~q ),
	.prn(vcc));
defparam \mem_used[70] .is_wysiwyg = "true";
defparam \mem_used[70] .power_up = "low";

cycloneive_lcell_comb \mem_used~120 (
	.dataa(\mem_used[68]~q ),
	.datab(\mem_used[70]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~120_combout ),
	.cout());
defparam \mem_used~120 .lut_mask = 16'hAACC;
defparam \mem_used~120 .sum_lutc_input = "datac";

dffeas \mem_used[69] (
	.clk(clk),
	.d(\mem_used~120_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[69]~q ),
	.prn(vcc));
defparam \mem_used[69] .is_wysiwyg = "true";
defparam \mem_used[69] .power_up = "low";

cycloneive_lcell_comb \mem_used~122 (
	.dataa(\mem_used[67]~q ),
	.datab(\mem_used[69]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~122_combout ),
	.cout());
defparam \mem_used~122 .lut_mask = 16'hAACC;
defparam \mem_used~122 .sum_lutc_input = "datac";

dffeas \mem_used[68] (
	.clk(clk),
	.d(\mem_used~122_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[68]~q ),
	.prn(vcc));
defparam \mem_used[68] .is_wysiwyg = "true";
defparam \mem_used[68] .power_up = "low";

cycloneive_lcell_comb \mem_used~124 (
	.dataa(\mem_used[66]~q ),
	.datab(\mem_used[68]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~124_combout ),
	.cout());
defparam \mem_used~124 .lut_mask = 16'hAACC;
defparam \mem_used~124 .sum_lutc_input = "datac";

dffeas \mem_used[67] (
	.clk(clk),
	.d(\mem_used~124_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[67]~q ),
	.prn(vcc));
defparam \mem_used[67] .is_wysiwyg = "true";
defparam \mem_used[67] .power_up = "low";

cycloneive_lcell_comb \mem_used~126 (
	.dataa(\mem_used[65]~q ),
	.datab(\mem_used[67]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~126_combout ),
	.cout());
defparam \mem_used~126 .lut_mask = 16'hAACC;
defparam \mem_used~126 .sum_lutc_input = "datac";

dffeas \mem_used[66] (
	.clk(clk),
	.d(\mem_used~126_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[66]~q ),
	.prn(vcc));
defparam \mem_used[66] .is_wysiwyg = "true";
defparam \mem_used[66] .power_up = "low";

cycloneive_lcell_comb \mem_used~128 (
	.dataa(\mem_used[64]~q ),
	.datab(\mem_used[66]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~128_combout ),
	.cout());
defparam \mem_used~128 .lut_mask = 16'hAACC;
defparam \mem_used~128 .sum_lutc_input = "datac";

dffeas \mem_used[65] (
	.clk(clk),
	.d(\mem_used~128_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[65]~q ),
	.prn(vcc));
defparam \mem_used[65] .is_wysiwyg = "true";
defparam \mem_used[65] .power_up = "low";

cycloneive_lcell_comb \mem_used~129 (
	.dataa(\mem_used[63]~q ),
	.datab(\mem_used[65]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~129_combout ),
	.cout());
defparam \mem_used~129 .lut_mask = 16'hAACC;
defparam \mem_used~129 .sum_lutc_input = "datac";

dffeas \mem_used[64] (
	.clk(clk),
	.d(\mem_used~129_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[64]~q ),
	.prn(vcc));
defparam \mem_used[64] .is_wysiwyg = "true";
defparam \mem_used[64] .power_up = "low";

cycloneive_lcell_comb \mem_used~127 (
	.dataa(\mem_used[62]~q ),
	.datab(\mem_used[64]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~127_combout ),
	.cout());
defparam \mem_used~127 .lut_mask = 16'hAACC;
defparam \mem_used~127 .sum_lutc_input = "datac";

dffeas \mem_used[63] (
	.clk(clk),
	.d(\mem_used~127_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[63]~q ),
	.prn(vcc));
defparam \mem_used[63] .is_wysiwyg = "true";
defparam \mem_used[63] .power_up = "low";

cycloneive_lcell_comb \mem_used~125 (
	.dataa(\mem_used[61]~q ),
	.datab(\mem_used[63]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~125_combout ),
	.cout());
defparam \mem_used~125 .lut_mask = 16'hAACC;
defparam \mem_used~125 .sum_lutc_input = "datac";

dffeas \mem_used[62] (
	.clk(clk),
	.d(\mem_used~125_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[62]~q ),
	.prn(vcc));
defparam \mem_used[62] .is_wysiwyg = "true";
defparam \mem_used[62] .power_up = "low";

cycloneive_lcell_comb \mem_used~123 (
	.dataa(\mem_used[60]~q ),
	.datab(\mem_used[62]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~123_combout ),
	.cout());
defparam \mem_used~123 .lut_mask = 16'hAACC;
defparam \mem_used~123 .sum_lutc_input = "datac";

dffeas \mem_used[61] (
	.clk(clk),
	.d(\mem_used~123_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[61]~q ),
	.prn(vcc));
defparam \mem_used[61] .is_wysiwyg = "true";
defparam \mem_used[61] .power_up = "low";

cycloneive_lcell_comb \mem_used~121 (
	.dataa(\mem_used[59]~q ),
	.datab(\mem_used[61]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~121_combout ),
	.cout());
defparam \mem_used~121 .lut_mask = 16'hAACC;
defparam \mem_used~121 .sum_lutc_input = "datac";

dffeas \mem_used[60] (
	.clk(clk),
	.d(\mem_used~121_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[60]~q ),
	.prn(vcc));
defparam \mem_used[60] .is_wysiwyg = "true";
defparam \mem_used[60] .power_up = "low";

cycloneive_lcell_comb \mem_used~119 (
	.dataa(\mem_used[58]~q ),
	.datab(\mem_used[60]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~119_combout ),
	.cout());
defparam \mem_used~119 .lut_mask = 16'hAACC;
defparam \mem_used~119 .sum_lutc_input = "datac";

dffeas \mem_used[59] (
	.clk(clk),
	.d(\mem_used~119_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[59]~q ),
	.prn(vcc));
defparam \mem_used[59] .is_wysiwyg = "true";
defparam \mem_used[59] .power_up = "low";

cycloneive_lcell_comb \mem_used~117 (
	.dataa(\mem_used[57]~q ),
	.datab(\mem_used[59]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~117_combout ),
	.cout());
defparam \mem_used~117 .lut_mask = 16'hAACC;
defparam \mem_used~117 .sum_lutc_input = "datac";

dffeas \mem_used[58] (
	.clk(clk),
	.d(\mem_used~117_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[58]~q ),
	.prn(vcc));
defparam \mem_used[58] .is_wysiwyg = "true";
defparam \mem_used[58] .power_up = "low";

cycloneive_lcell_comb \mem_used~115 (
	.dataa(\mem_used[56]~q ),
	.datab(\mem_used[58]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~115_combout ),
	.cout());
defparam \mem_used~115 .lut_mask = 16'hAACC;
defparam \mem_used~115 .sum_lutc_input = "datac";

dffeas \mem_used[57] (
	.clk(clk),
	.d(\mem_used~115_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[57]~q ),
	.prn(vcc));
defparam \mem_used[57] .is_wysiwyg = "true";
defparam \mem_used[57] .power_up = "low";

cycloneive_lcell_comb \mem_used~113 (
	.dataa(\mem_used[55]~q ),
	.datab(\mem_used[57]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~113_combout ),
	.cout());
defparam \mem_used~113 .lut_mask = 16'hAACC;
defparam \mem_used~113 .sum_lutc_input = "datac";

dffeas \mem_used[56] (
	.clk(clk),
	.d(\mem_used~113_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[56]~q ),
	.prn(vcc));
defparam \mem_used[56] .is_wysiwyg = "true";
defparam \mem_used[56] .power_up = "low";

cycloneive_lcell_comb \mem_used~111 (
	.dataa(\mem_used[54]~q ),
	.datab(\mem_used[56]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~111_combout ),
	.cout());
defparam \mem_used~111 .lut_mask = 16'hAACC;
defparam \mem_used~111 .sum_lutc_input = "datac";

dffeas \mem_used[55] (
	.clk(clk),
	.d(\mem_used~111_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[55]~q ),
	.prn(vcc));
defparam \mem_used[55] .is_wysiwyg = "true";
defparam \mem_used[55] .power_up = "low";

cycloneive_lcell_comb \mem_used~109 (
	.dataa(\mem_used[53]~q ),
	.datab(\mem_used[55]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~109_combout ),
	.cout());
defparam \mem_used~109 .lut_mask = 16'hAACC;
defparam \mem_used~109 .sum_lutc_input = "datac";

dffeas \mem_used[54] (
	.clk(clk),
	.d(\mem_used~109_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[54]~q ),
	.prn(vcc));
defparam \mem_used[54] .is_wysiwyg = "true";
defparam \mem_used[54] .power_up = "low";

cycloneive_lcell_comb \mem_used~107 (
	.dataa(\mem_used[52]~q ),
	.datab(\mem_used[54]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~107_combout ),
	.cout());
defparam \mem_used~107 .lut_mask = 16'hAACC;
defparam \mem_used~107 .sum_lutc_input = "datac";

dffeas \mem_used[53] (
	.clk(clk),
	.d(\mem_used~107_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[53]~q ),
	.prn(vcc));
defparam \mem_used[53] .is_wysiwyg = "true";
defparam \mem_used[53] .power_up = "low";

cycloneive_lcell_comb \mem_used~105 (
	.dataa(\mem_used[51]~q ),
	.datab(\mem_used[53]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~105_combout ),
	.cout());
defparam \mem_used~105 .lut_mask = 16'hAACC;
defparam \mem_used~105 .sum_lutc_input = "datac";

dffeas \mem_used[52] (
	.clk(clk),
	.d(\mem_used~105_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[52]~q ),
	.prn(vcc));
defparam \mem_used[52] .is_wysiwyg = "true";
defparam \mem_used[52] .power_up = "low";

cycloneive_lcell_comb \mem_used~103 (
	.dataa(\mem_used[50]~q ),
	.datab(\mem_used[52]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~103_combout ),
	.cout());
defparam \mem_used~103 .lut_mask = 16'hAACC;
defparam \mem_used~103 .sum_lutc_input = "datac";

dffeas \mem_used[51] (
	.clk(clk),
	.d(\mem_used~103_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[51]~q ),
	.prn(vcc));
defparam \mem_used[51] .is_wysiwyg = "true";
defparam \mem_used[51] .power_up = "low";

cycloneive_lcell_comb \mem_used~101 (
	.dataa(\mem_used[49]~q ),
	.datab(\mem_used[51]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~101_combout ),
	.cout());
defparam \mem_used~101 .lut_mask = 16'hAACC;
defparam \mem_used~101 .sum_lutc_input = "datac";

dffeas \mem_used[50] (
	.clk(clk),
	.d(\mem_used~101_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[50]~q ),
	.prn(vcc));
defparam \mem_used[50] .is_wysiwyg = "true";
defparam \mem_used[50] .power_up = "low";

cycloneive_lcell_comb \mem_used~99 (
	.dataa(\mem_used[48]~q ),
	.datab(\mem_used[50]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~99_combout ),
	.cout());
defparam \mem_used~99 .lut_mask = 16'hAACC;
defparam \mem_used~99 .sum_lutc_input = "datac";

dffeas \mem_used[49] (
	.clk(clk),
	.d(\mem_used~99_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[49]~q ),
	.prn(vcc));
defparam \mem_used[49] .is_wysiwyg = "true";
defparam \mem_used[49] .power_up = "low";

cycloneive_lcell_comb \mem_used~97 (
	.dataa(\mem_used[47]~q ),
	.datab(\mem_used[49]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~97_combout ),
	.cout());
defparam \mem_used~97 .lut_mask = 16'hAACC;
defparam \mem_used~97 .sum_lutc_input = "datac";

dffeas \mem_used[48] (
	.clk(clk),
	.d(\mem_used~97_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[48]~q ),
	.prn(vcc));
defparam \mem_used[48] .is_wysiwyg = "true";
defparam \mem_used[48] .power_up = "low";

cycloneive_lcell_comb \mem_used~95 (
	.dataa(\mem_used[46]~q ),
	.datab(\mem_used[48]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~95_combout ),
	.cout());
defparam \mem_used~95 .lut_mask = 16'hAACC;
defparam \mem_used~95 .sum_lutc_input = "datac";

dffeas \mem_used[47] (
	.clk(clk),
	.d(\mem_used~95_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[47]~q ),
	.prn(vcc));
defparam \mem_used[47] .is_wysiwyg = "true";
defparam \mem_used[47] .power_up = "low";

cycloneive_lcell_comb \mem_used~93 (
	.dataa(\mem_used[45]~q ),
	.datab(\mem_used[47]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~93_combout ),
	.cout());
defparam \mem_used~93 .lut_mask = 16'hAACC;
defparam \mem_used~93 .sum_lutc_input = "datac";

dffeas \mem_used[46] (
	.clk(clk),
	.d(\mem_used~93_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[46]~q ),
	.prn(vcc));
defparam \mem_used[46] .is_wysiwyg = "true";
defparam \mem_used[46] .power_up = "low";

cycloneive_lcell_comb \mem_used~91 (
	.dataa(\mem_used[44]~q ),
	.datab(\mem_used[46]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~91_combout ),
	.cout());
defparam \mem_used~91 .lut_mask = 16'hAACC;
defparam \mem_used~91 .sum_lutc_input = "datac";

dffeas \mem_used[45] (
	.clk(clk),
	.d(\mem_used~91_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[45]~q ),
	.prn(vcc));
defparam \mem_used[45] .is_wysiwyg = "true";
defparam \mem_used[45] .power_up = "low";

cycloneive_lcell_comb \mem_used~89 (
	.dataa(\mem_used[43]~q ),
	.datab(\mem_used[45]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~89_combout ),
	.cout());
defparam \mem_used~89 .lut_mask = 16'hAACC;
defparam \mem_used~89 .sum_lutc_input = "datac";

dffeas \mem_used[44] (
	.clk(clk),
	.d(\mem_used~89_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[44]~q ),
	.prn(vcc));
defparam \mem_used[44] .is_wysiwyg = "true";
defparam \mem_used[44] .power_up = "low";

cycloneive_lcell_comb \mem_used~87 (
	.dataa(\mem_used[42]~q ),
	.datab(\mem_used[44]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~87_combout ),
	.cout());
defparam \mem_used~87 .lut_mask = 16'hAACC;
defparam \mem_used~87 .sum_lutc_input = "datac";

dffeas \mem_used[43] (
	.clk(clk),
	.d(\mem_used~87_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[43]~q ),
	.prn(vcc));
defparam \mem_used[43] .is_wysiwyg = "true";
defparam \mem_used[43] .power_up = "low";

cycloneive_lcell_comb \mem_used~85 (
	.dataa(\mem_used[41]~q ),
	.datab(\mem_used[43]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~85_combout ),
	.cout());
defparam \mem_used~85 .lut_mask = 16'hAACC;
defparam \mem_used~85 .sum_lutc_input = "datac";

dffeas \mem_used[42] (
	.clk(clk),
	.d(\mem_used~85_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[42]~q ),
	.prn(vcc));
defparam \mem_used[42] .is_wysiwyg = "true";
defparam \mem_used[42] .power_up = "low";

cycloneive_lcell_comb \mem_used~83 (
	.dataa(\mem_used[40]~q ),
	.datab(\mem_used[42]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~83_combout ),
	.cout());
defparam \mem_used~83 .lut_mask = 16'hAACC;
defparam \mem_used~83 .sum_lutc_input = "datac";

dffeas \mem_used[41] (
	.clk(clk),
	.d(\mem_used~83_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[41]~q ),
	.prn(vcc));
defparam \mem_used[41] .is_wysiwyg = "true";
defparam \mem_used[41] .power_up = "low";

cycloneive_lcell_comb \mem_used~81 (
	.dataa(\mem_used[39]~q ),
	.datab(\mem_used[41]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~81_combout ),
	.cout());
defparam \mem_used~81 .lut_mask = 16'hAACC;
defparam \mem_used~81 .sum_lutc_input = "datac";

dffeas \mem_used[40] (
	.clk(clk),
	.d(\mem_used~81_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[40]~q ),
	.prn(vcc));
defparam \mem_used[40] .is_wysiwyg = "true";
defparam \mem_used[40] .power_up = "low";

cycloneive_lcell_comb \mem_used~79 (
	.dataa(\mem_used[38]~q ),
	.datab(\mem_used[40]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~79_combout ),
	.cout());
defparam \mem_used~79 .lut_mask = 16'hAACC;
defparam \mem_used~79 .sum_lutc_input = "datac";

dffeas \mem_used[39] (
	.clk(clk),
	.d(\mem_used~79_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[39]~q ),
	.prn(vcc));
defparam \mem_used[39] .is_wysiwyg = "true";
defparam \mem_used[39] .power_up = "low";

cycloneive_lcell_comb \mem_used~77 (
	.dataa(\mem_used[37]~q ),
	.datab(\mem_used[39]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~77_combout ),
	.cout());
defparam \mem_used~77 .lut_mask = 16'hAACC;
defparam \mem_used~77 .sum_lutc_input = "datac";

dffeas \mem_used[38] (
	.clk(clk),
	.d(\mem_used~77_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[38]~q ),
	.prn(vcc));
defparam \mem_used[38] .is_wysiwyg = "true";
defparam \mem_used[38] .power_up = "low";

cycloneive_lcell_comb \mem_used~75 (
	.dataa(\mem_used[36]~q ),
	.datab(\mem_used[38]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~75_combout ),
	.cout());
defparam \mem_used~75 .lut_mask = 16'hAACC;
defparam \mem_used~75 .sum_lutc_input = "datac";

dffeas \mem_used[37] (
	.clk(clk),
	.d(\mem_used~75_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[37]~q ),
	.prn(vcc));
defparam \mem_used[37] .is_wysiwyg = "true";
defparam \mem_used[37] .power_up = "low";

cycloneive_lcell_comb \mem_used~73 (
	.dataa(\mem_used[35]~q ),
	.datab(\mem_used[37]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~73_combout ),
	.cout());
defparam \mem_used~73 .lut_mask = 16'hAACC;
defparam \mem_used~73 .sum_lutc_input = "datac";

dffeas \mem_used[36] (
	.clk(clk),
	.d(\mem_used~73_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[36]~q ),
	.prn(vcc));
defparam \mem_used[36] .is_wysiwyg = "true";
defparam \mem_used[36] .power_up = "low";

cycloneive_lcell_comb \mem_used~71 (
	.dataa(\mem_used[34]~q ),
	.datab(\mem_used[36]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~71_combout ),
	.cout());
defparam \mem_used~71 .lut_mask = 16'hAACC;
defparam \mem_used~71 .sum_lutc_input = "datac";

dffeas \mem_used[35] (
	.clk(clk),
	.d(\mem_used~71_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[35]~q ),
	.prn(vcc));
defparam \mem_used[35] .is_wysiwyg = "true";
defparam \mem_used[35] .power_up = "low";

cycloneive_lcell_comb \mem_used~69 (
	.dataa(\mem_used[33]~q ),
	.datab(\mem_used[35]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~69_combout ),
	.cout());
defparam \mem_used~69 .lut_mask = 16'hAACC;
defparam \mem_used~69 .sum_lutc_input = "datac";

dffeas \mem_used[34] (
	.clk(clk),
	.d(\mem_used~69_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[34]~q ),
	.prn(vcc));
defparam \mem_used[34] .is_wysiwyg = "true";
defparam \mem_used[34] .power_up = "low";

cycloneive_lcell_comb \mem_used~67 (
	.dataa(\mem_used[32]~q ),
	.datab(\mem_used[34]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~67_combout ),
	.cout());
defparam \mem_used~67 .lut_mask = 16'hAACC;
defparam \mem_used~67 .sum_lutc_input = "datac";

dffeas \mem_used[33] (
	.clk(clk),
	.d(\mem_used~67_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[33]~q ),
	.prn(vcc));
defparam \mem_used[33] .is_wysiwyg = "true";
defparam \mem_used[33] .power_up = "low";

cycloneive_lcell_comb \mem_used~65 (
	.dataa(\mem_used[31]~q ),
	.datab(\mem_used[33]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~65_combout ),
	.cout());
defparam \mem_used~65 .lut_mask = 16'hAACC;
defparam \mem_used~65 .sum_lutc_input = "datac";

dffeas \mem_used[32] (
	.clk(clk),
	.d(\mem_used~65_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[32]~q ),
	.prn(vcc));
defparam \mem_used[32] .is_wysiwyg = "true";
defparam \mem_used[32] .power_up = "low";

cycloneive_lcell_comb \mem_used~63 (
	.dataa(\mem_used[30]~q ),
	.datab(\mem_used[32]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~63_combout ),
	.cout());
defparam \mem_used~63 .lut_mask = 16'hAACC;
defparam \mem_used~63 .sum_lutc_input = "datac";

dffeas \mem_used[31] (
	.clk(clk),
	.d(\mem_used~63_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[31]~q ),
	.prn(vcc));
defparam \mem_used[31] .is_wysiwyg = "true";
defparam \mem_used[31] .power_up = "low";

cycloneive_lcell_comb \mem_used~61 (
	.dataa(\mem_used[29]~q ),
	.datab(\mem_used[31]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~61_combout ),
	.cout());
defparam \mem_used~61 .lut_mask = 16'hAACC;
defparam \mem_used~61 .sum_lutc_input = "datac";

dffeas \mem_used[30] (
	.clk(clk),
	.d(\mem_used~61_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[30]~q ),
	.prn(vcc));
defparam \mem_used[30] .is_wysiwyg = "true";
defparam \mem_used[30] .power_up = "low";

cycloneive_lcell_comb \mem_used~59 (
	.dataa(\mem_used[28]~q ),
	.datab(\mem_used[30]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~59_combout ),
	.cout());
defparam \mem_used~59 .lut_mask = 16'hAACC;
defparam \mem_used~59 .sum_lutc_input = "datac";

dffeas \mem_used[29] (
	.clk(clk),
	.d(\mem_used~59_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[29]~q ),
	.prn(vcc));
defparam \mem_used[29] .is_wysiwyg = "true";
defparam \mem_used[29] .power_up = "low";

cycloneive_lcell_comb \mem_used~57 (
	.dataa(\mem_used[27]~q ),
	.datab(\mem_used[29]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~57_combout ),
	.cout());
defparam \mem_used~57 .lut_mask = 16'hAACC;
defparam \mem_used~57 .sum_lutc_input = "datac";

dffeas \mem_used[28] (
	.clk(clk),
	.d(\mem_used~57_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[28]~q ),
	.prn(vcc));
defparam \mem_used[28] .is_wysiwyg = "true";
defparam \mem_used[28] .power_up = "low";

cycloneive_lcell_comb \mem_used~55 (
	.dataa(\mem_used[26]~q ),
	.datab(\mem_used[28]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~55_combout ),
	.cout());
defparam \mem_used~55 .lut_mask = 16'hAACC;
defparam \mem_used~55 .sum_lutc_input = "datac";

dffeas \mem_used[27] (
	.clk(clk),
	.d(\mem_used~55_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[27]~q ),
	.prn(vcc));
defparam \mem_used[27] .is_wysiwyg = "true";
defparam \mem_used[27] .power_up = "low";

cycloneive_lcell_comb \mem_used~53 (
	.dataa(\mem_used[25]~q ),
	.datab(\mem_used[27]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~53_combout ),
	.cout());
defparam \mem_used~53 .lut_mask = 16'hAACC;
defparam \mem_used~53 .sum_lutc_input = "datac";

dffeas \mem_used[26] (
	.clk(clk),
	.d(\mem_used~53_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[26]~q ),
	.prn(vcc));
defparam \mem_used[26] .is_wysiwyg = "true";
defparam \mem_used[26] .power_up = "low";

cycloneive_lcell_comb \mem_used~51 (
	.dataa(\mem_used[24]~q ),
	.datab(\mem_used[26]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~51_combout ),
	.cout());
defparam \mem_used~51 .lut_mask = 16'hAACC;
defparam \mem_used~51 .sum_lutc_input = "datac";

dffeas \mem_used[25] (
	.clk(clk),
	.d(\mem_used~51_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[25]~q ),
	.prn(vcc));
defparam \mem_used[25] .is_wysiwyg = "true";
defparam \mem_used[25] .power_up = "low";

cycloneive_lcell_comb \mem_used~49 (
	.dataa(\mem_used[23]~q ),
	.datab(\mem_used[25]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~49_combout ),
	.cout());
defparam \mem_used~49 .lut_mask = 16'hAACC;
defparam \mem_used~49 .sum_lutc_input = "datac";

dffeas \mem_used[24] (
	.clk(clk),
	.d(\mem_used~49_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[24]~q ),
	.prn(vcc));
defparam \mem_used[24] .is_wysiwyg = "true";
defparam \mem_used[24] .power_up = "low";

cycloneive_lcell_comb \mem_used~47 (
	.dataa(\mem_used[22]~q ),
	.datab(\mem_used[24]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~47_combout ),
	.cout());
defparam \mem_used~47 .lut_mask = 16'hAACC;
defparam \mem_used~47 .sum_lutc_input = "datac";

dffeas \mem_used[23] (
	.clk(clk),
	.d(\mem_used~47_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[23]~q ),
	.prn(vcc));
defparam \mem_used[23] .is_wysiwyg = "true";
defparam \mem_used[23] .power_up = "low";

cycloneive_lcell_comb \mem_used~45 (
	.dataa(\mem_used[21]~q ),
	.datab(\mem_used[23]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~45_combout ),
	.cout());
defparam \mem_used~45 .lut_mask = 16'hAACC;
defparam \mem_used~45 .sum_lutc_input = "datac";

dffeas \mem_used[22] (
	.clk(clk),
	.d(\mem_used~45_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[22]~q ),
	.prn(vcc));
defparam \mem_used[22] .is_wysiwyg = "true";
defparam \mem_used[22] .power_up = "low";

cycloneive_lcell_comb \mem_used~43 (
	.dataa(\mem_used[20]~q ),
	.datab(\mem_used[22]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~43_combout ),
	.cout());
defparam \mem_used~43 .lut_mask = 16'hAACC;
defparam \mem_used~43 .sum_lutc_input = "datac";

dffeas \mem_used[21] (
	.clk(clk),
	.d(\mem_used~43_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[21]~q ),
	.prn(vcc));
defparam \mem_used[21] .is_wysiwyg = "true";
defparam \mem_used[21] .power_up = "low";

cycloneive_lcell_comb \mem_used~41 (
	.dataa(\mem_used[19]~q ),
	.datab(\mem_used[21]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~41_combout ),
	.cout());
defparam \mem_used~41 .lut_mask = 16'hAACC;
defparam \mem_used~41 .sum_lutc_input = "datac";

dffeas \mem_used[20] (
	.clk(clk),
	.d(\mem_used~41_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[20]~q ),
	.prn(vcc));
defparam \mem_used[20] .is_wysiwyg = "true";
defparam \mem_used[20] .power_up = "low";

cycloneive_lcell_comb \mem_used~39 (
	.dataa(\mem_used[18]~q ),
	.datab(\mem_used[20]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~39_combout ),
	.cout());
defparam \mem_used~39 .lut_mask = 16'hAACC;
defparam \mem_used~39 .sum_lutc_input = "datac";

dffeas \mem_used[19] (
	.clk(clk),
	.d(\mem_used~39_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[19]~q ),
	.prn(vcc));
defparam \mem_used[19] .is_wysiwyg = "true";
defparam \mem_used[19] .power_up = "low";

cycloneive_lcell_comb \mem_used~37 (
	.dataa(\mem_used[17]~q ),
	.datab(\mem_used[19]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~37_combout ),
	.cout());
defparam \mem_used~37 .lut_mask = 16'hAACC;
defparam \mem_used~37 .sum_lutc_input = "datac";

dffeas \mem_used[18] (
	.clk(clk),
	.d(\mem_used~37_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[18]~q ),
	.prn(vcc));
defparam \mem_used[18] .is_wysiwyg = "true";
defparam \mem_used[18] .power_up = "low";

cycloneive_lcell_comb \mem_used~35 (
	.dataa(\mem_used[16]~q ),
	.datab(\mem_used[18]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~35_combout ),
	.cout());
defparam \mem_used~35 .lut_mask = 16'hAACC;
defparam \mem_used~35 .sum_lutc_input = "datac";

dffeas \mem_used[17] (
	.clk(clk),
	.d(\mem_used~35_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[17]~q ),
	.prn(vcc));
defparam \mem_used[17] .is_wysiwyg = "true";
defparam \mem_used[17] .power_up = "low";

cycloneive_lcell_comb \mem_used~33 (
	.dataa(\mem_used[15]~q ),
	.datab(\mem_used[17]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~33_combout ),
	.cout());
defparam \mem_used~33 .lut_mask = 16'hAACC;
defparam \mem_used~33 .sum_lutc_input = "datac";

dffeas \mem_used[16] (
	.clk(clk),
	.d(\mem_used~33_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[16]~q ),
	.prn(vcc));
defparam \mem_used[16] .is_wysiwyg = "true";
defparam \mem_used[16] .power_up = "low";

cycloneive_lcell_comb \mem_used~31 (
	.dataa(\mem_used[14]~q ),
	.datab(\mem_used[16]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~31_combout ),
	.cout());
defparam \mem_used~31 .lut_mask = 16'hAACC;
defparam \mem_used~31 .sum_lutc_input = "datac";

dffeas \mem_used[15] (
	.clk(clk),
	.d(\mem_used~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[15]~q ),
	.prn(vcc));
defparam \mem_used[15] .is_wysiwyg = "true";
defparam \mem_used[15] .power_up = "low";

cycloneive_lcell_comb \mem_used~29 (
	.dataa(\mem_used[13]~q ),
	.datab(\mem_used[15]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~29_combout ),
	.cout());
defparam \mem_used~29 .lut_mask = 16'hAACC;
defparam \mem_used~29 .sum_lutc_input = "datac";

dffeas \mem_used[14] (
	.clk(clk),
	.d(\mem_used~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[14]~q ),
	.prn(vcc));
defparam \mem_used[14] .is_wysiwyg = "true";
defparam \mem_used[14] .power_up = "low";

cycloneive_lcell_comb \mem_used~27 (
	.dataa(\mem_used[12]~q ),
	.datab(\mem_used[14]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~27_combout ),
	.cout());
defparam \mem_used~27 .lut_mask = 16'hAACC;
defparam \mem_used~27 .sum_lutc_input = "datac";

dffeas \mem_used[13] (
	.clk(clk),
	.d(\mem_used~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[13]~q ),
	.prn(vcc));
defparam \mem_used[13] .is_wysiwyg = "true";
defparam \mem_used[13] .power_up = "low";

cycloneive_lcell_comb \mem_used~25 (
	.dataa(\mem_used[11]~q ),
	.datab(\mem_used[13]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~25_combout ),
	.cout());
defparam \mem_used~25 .lut_mask = 16'hAACC;
defparam \mem_used~25 .sum_lutc_input = "datac";

dffeas \mem_used[12] (
	.clk(clk),
	.d(\mem_used~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[12]~q ),
	.prn(vcc));
defparam \mem_used[12] .is_wysiwyg = "true";
defparam \mem_used[12] .power_up = "low";

cycloneive_lcell_comb \mem_used~23 (
	.dataa(\mem_used[10]~q ),
	.datab(\mem_used[12]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~23_combout ),
	.cout());
defparam \mem_used~23 .lut_mask = 16'hAACC;
defparam \mem_used~23 .sum_lutc_input = "datac";

dffeas \mem_used[11] (
	.clk(clk),
	.d(\mem_used~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[11]~q ),
	.prn(vcc));
defparam \mem_used[11] .is_wysiwyg = "true";
defparam \mem_used[11] .power_up = "low";

cycloneive_lcell_comb \mem_used~21 (
	.dataa(\mem_used[9]~q ),
	.datab(\mem_used[11]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~21_combout ),
	.cout());
defparam \mem_used~21 .lut_mask = 16'hAACC;
defparam \mem_used~21 .sum_lutc_input = "datac";

dffeas \mem_used[10] (
	.clk(clk),
	.d(\mem_used~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[10]~q ),
	.prn(vcc));
defparam \mem_used[10] .is_wysiwyg = "true";
defparam \mem_used[10] .power_up = "low";

cycloneive_lcell_comb \mem_used~19 (
	.dataa(\mem_used[8]~q ),
	.datab(\mem_used[10]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~19_combout ),
	.cout());
defparam \mem_used~19 .lut_mask = 16'hAACC;
defparam \mem_used~19 .sum_lutc_input = "datac";

dffeas \mem_used[9] (
	.clk(clk),
	.d(\mem_used~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[9]~q ),
	.prn(vcc));
defparam \mem_used[9] .is_wysiwyg = "true";
defparam \mem_used[9] .power_up = "low";

cycloneive_lcell_comb \mem_used~17 (
	.dataa(\mem_used[7]~q ),
	.datab(\mem_used[9]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~17_combout ),
	.cout());
defparam \mem_used~17 .lut_mask = 16'hAACC;
defparam \mem_used~17 .sum_lutc_input = "datac";

dffeas \mem_used[8] (
	.clk(clk),
	.d(\mem_used~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[8]~q ),
	.prn(vcc));
defparam \mem_used[8] .is_wysiwyg = "true";
defparam \mem_used[8] .power_up = "low";

cycloneive_lcell_comb \mem_used~15 (
	.dataa(\mem_used[6]~q ),
	.datab(\mem_used[8]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~15_combout ),
	.cout());
defparam \mem_used~15 .lut_mask = 16'hAACC;
defparam \mem_used~15 .sum_lutc_input = "datac";

dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[7]~q ),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

cycloneive_lcell_comb \mem_used~13 (
	.dataa(\mem_used[5]~q ),
	.datab(\mem_used[7]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~13_combout ),
	.cout());
defparam \mem_used~13 .lut_mask = 16'hAACC;
defparam \mem_used~13 .sum_lutc_input = "datac";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cycloneive_lcell_comb \mem_used~11 (
	.dataa(\mem_used[4]~q ),
	.datab(\mem_used[6]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~11_combout ),
	.cout());
defparam \mem_used~11 .lut_mask = 16'hAACC;
defparam \mem_used~11 .sum_lutc_input = "datac";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cycloneive_lcell_comb \mem_used~9 (
	.dataa(\mem_used[3]~q ),
	.datab(\mem_used[5]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~9_combout ),
	.cout());
defparam \mem_used~9 .lut_mask = 16'hAACC;
defparam \mem_used~9 .sum_lutc_input = "datac";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cycloneive_lcell_comb \mem_used~7 (
	.dataa(\mem_used[2]~q ),
	.datab(\mem_used[4]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~7_combout ),
	.cout());
defparam \mem_used~7 .lut_mask = 16'hAACC;
defparam \mem_used~7 .sum_lutc_input = "datac";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cycloneive_lcell_comb \mem_used~5 (
	.dataa(\mem_used[1]~q ),
	.datab(\mem_used[3]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~5_combout ),
	.cout());
defparam \mem_used~5 .lut_mask = 16'hAACC;
defparam \mem_used~5 .sum_lutc_input = "datac";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cycloneive_lcell_comb \mem_used~1 (
	.dataa(\mem_used[0]~q ),
	.datab(\mem_used[2]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~1_combout ),
	.cout());
defparam \mem_used~1 .lut_mask = 16'hAACC;
defparam \mem_used~1 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[127]~2_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\write~0_combout ),
	.datab(\mem_used[0]~q ),
	.datac(\mem_used[1]~q ),
	.datad(out_valid),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \read~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(out_valid),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h0FFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[127][67]~255 (
	.dataa(\mem[127][67]~q ),
	.datab(\mem~254_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[127]~q ),
	.cin(gnd),
	.combout(\mem[127][67]~255_combout ),
	.cout());
defparam \mem[127][67]~255 .lut_mask = 16'hEFFE;
defparam \mem[127][67]~255 .sum_lutc_input = "datac";

dffeas \mem[127][67] (
	.clk(clk),
	.d(\mem[127][67]~255_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[127][67]~q ),
	.prn(vcc));
defparam \mem[127][67] .is_wysiwyg = "true";
defparam \mem[127][67] .power_up = "low";

cycloneive_lcell_comb \mem[126][67]~252 (
	.dataa(\mem[127][67]~q ),
	.datab(\mem_used[127]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[126][67]~252_combout ),
	.cout());
defparam \mem[126][67]~252 .lut_mask = 16'hB8FF;
defparam \mem[126][67]~252 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[126][67]~253 (
	.dataa(\mem[126][67]~q ),
	.datab(\mem[126][67]~252_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[126]~q ),
	.cin(gnd),
	.combout(\mem[126][67]~253_combout ),
	.cout());
defparam \mem[126][67]~253 .lut_mask = 16'hEFFE;
defparam \mem[126][67]~253 .sum_lutc_input = "datac";

dffeas \mem[126][67] (
	.clk(clk),
	.d(\mem[126][67]~253_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[126][67]~q ),
	.prn(vcc));
defparam \mem[126][67] .is_wysiwyg = "true";
defparam \mem[126][67] .power_up = "low";

cycloneive_lcell_comb \mem[125][67]~250 (
	.dataa(\mem[126][67]~q ),
	.datab(\mem_used[126]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[125][67]~250_combout ),
	.cout());
defparam \mem[125][67]~250 .lut_mask = 16'hB8FF;
defparam \mem[125][67]~250 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[125][67]~251 (
	.dataa(\mem[125][67]~q ),
	.datab(\mem[125][67]~250_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[125]~q ),
	.cin(gnd),
	.combout(\mem[125][67]~251_combout ),
	.cout());
defparam \mem[125][67]~251 .lut_mask = 16'hEFFE;
defparam \mem[125][67]~251 .sum_lutc_input = "datac";

dffeas \mem[125][67] (
	.clk(clk),
	.d(\mem[125][67]~251_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[125][67]~q ),
	.prn(vcc));
defparam \mem[125][67] .is_wysiwyg = "true";
defparam \mem[125][67] .power_up = "low";

cycloneive_lcell_comb \mem[124][67]~248 (
	.dataa(\mem[125][67]~q ),
	.datab(\mem_used[125]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[124][67]~248_combout ),
	.cout());
defparam \mem[124][67]~248 .lut_mask = 16'hB8FF;
defparam \mem[124][67]~248 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[124][67]~249 (
	.dataa(\mem[124][67]~q ),
	.datab(\mem[124][67]~248_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[124]~q ),
	.cin(gnd),
	.combout(\mem[124][67]~249_combout ),
	.cout());
defparam \mem[124][67]~249 .lut_mask = 16'hEFFE;
defparam \mem[124][67]~249 .sum_lutc_input = "datac";

dffeas \mem[124][67] (
	.clk(clk),
	.d(\mem[124][67]~249_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[124][67]~q ),
	.prn(vcc));
defparam \mem[124][67] .is_wysiwyg = "true";
defparam \mem[124][67] .power_up = "low";

cycloneive_lcell_comb \mem[123][67]~246 (
	.dataa(\mem[124][67]~q ),
	.datab(\mem_used[124]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[123][67]~246_combout ),
	.cout());
defparam \mem[123][67]~246 .lut_mask = 16'hB8FF;
defparam \mem[123][67]~246 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[123][67]~247 (
	.dataa(\mem[123][67]~q ),
	.datab(\mem[123][67]~246_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[123]~q ),
	.cin(gnd),
	.combout(\mem[123][67]~247_combout ),
	.cout());
defparam \mem[123][67]~247 .lut_mask = 16'hEFFE;
defparam \mem[123][67]~247 .sum_lutc_input = "datac";

dffeas \mem[123][67] (
	.clk(clk),
	.d(\mem[123][67]~247_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[123][67]~q ),
	.prn(vcc));
defparam \mem[123][67] .is_wysiwyg = "true";
defparam \mem[123][67] .power_up = "low";

cycloneive_lcell_comb \mem[122][67]~244 (
	.dataa(\mem[123][67]~q ),
	.datab(\mem_used[123]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[122][67]~244_combout ),
	.cout());
defparam \mem[122][67]~244 .lut_mask = 16'hB8FF;
defparam \mem[122][67]~244 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[122][67]~245 (
	.dataa(\mem[122][67]~q ),
	.datab(\mem[122][67]~244_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[122]~q ),
	.cin(gnd),
	.combout(\mem[122][67]~245_combout ),
	.cout());
defparam \mem[122][67]~245 .lut_mask = 16'hEFFE;
defparam \mem[122][67]~245 .sum_lutc_input = "datac";

dffeas \mem[122][67] (
	.clk(clk),
	.d(\mem[122][67]~245_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[122][67]~q ),
	.prn(vcc));
defparam \mem[122][67] .is_wysiwyg = "true";
defparam \mem[122][67] .power_up = "low";

cycloneive_lcell_comb \mem[121][67]~242 (
	.dataa(\mem[122][67]~q ),
	.datab(\mem_used[122]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[121][67]~242_combout ),
	.cout());
defparam \mem[121][67]~242 .lut_mask = 16'hB8FF;
defparam \mem[121][67]~242 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[121][67]~243 (
	.dataa(\mem[121][67]~q ),
	.datab(\mem[121][67]~242_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[121]~q ),
	.cin(gnd),
	.combout(\mem[121][67]~243_combout ),
	.cout());
defparam \mem[121][67]~243 .lut_mask = 16'hEFFE;
defparam \mem[121][67]~243 .sum_lutc_input = "datac";

dffeas \mem[121][67] (
	.clk(clk),
	.d(\mem[121][67]~243_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[121][67]~q ),
	.prn(vcc));
defparam \mem[121][67] .is_wysiwyg = "true";
defparam \mem[121][67] .power_up = "low";

cycloneive_lcell_comb \mem[120][67]~240 (
	.dataa(\mem[121][67]~q ),
	.datab(\mem_used[121]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[120][67]~240_combout ),
	.cout());
defparam \mem[120][67]~240 .lut_mask = 16'hB8FF;
defparam \mem[120][67]~240 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[120][67]~241 (
	.dataa(\mem[120][67]~q ),
	.datab(\mem[120][67]~240_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[120]~q ),
	.cin(gnd),
	.combout(\mem[120][67]~241_combout ),
	.cout());
defparam \mem[120][67]~241 .lut_mask = 16'hEFFE;
defparam \mem[120][67]~241 .sum_lutc_input = "datac";

dffeas \mem[120][67] (
	.clk(clk),
	.d(\mem[120][67]~241_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[120][67]~q ),
	.prn(vcc));
defparam \mem[120][67] .is_wysiwyg = "true";
defparam \mem[120][67] .power_up = "low";

cycloneive_lcell_comb \mem[119][67]~238 (
	.dataa(\mem[120][67]~q ),
	.datab(\mem_used[120]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[119][67]~238_combout ),
	.cout());
defparam \mem[119][67]~238 .lut_mask = 16'hB8FF;
defparam \mem[119][67]~238 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[119][67]~239 (
	.dataa(\mem[119][67]~q ),
	.datab(\mem[119][67]~238_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[119]~q ),
	.cin(gnd),
	.combout(\mem[119][67]~239_combout ),
	.cout());
defparam \mem[119][67]~239 .lut_mask = 16'hEFFE;
defparam \mem[119][67]~239 .sum_lutc_input = "datac";

dffeas \mem[119][67] (
	.clk(clk),
	.d(\mem[119][67]~239_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[119][67]~q ),
	.prn(vcc));
defparam \mem[119][67] .is_wysiwyg = "true";
defparam \mem[119][67] .power_up = "low";

cycloneive_lcell_comb \mem[118][67]~236 (
	.dataa(\mem[119][67]~q ),
	.datab(\mem_used[119]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[118][67]~236_combout ),
	.cout());
defparam \mem[118][67]~236 .lut_mask = 16'hB8FF;
defparam \mem[118][67]~236 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[118][67]~237 (
	.dataa(\mem[118][67]~q ),
	.datab(\mem[118][67]~236_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[118]~q ),
	.cin(gnd),
	.combout(\mem[118][67]~237_combout ),
	.cout());
defparam \mem[118][67]~237 .lut_mask = 16'hEFFE;
defparam \mem[118][67]~237 .sum_lutc_input = "datac";

dffeas \mem[118][67] (
	.clk(clk),
	.d(\mem[118][67]~237_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[118][67]~q ),
	.prn(vcc));
defparam \mem[118][67] .is_wysiwyg = "true";
defparam \mem[118][67] .power_up = "low";

cycloneive_lcell_comb \mem[117][67]~234 (
	.dataa(\mem[118][67]~q ),
	.datab(\mem_used[118]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[117][67]~234_combout ),
	.cout());
defparam \mem[117][67]~234 .lut_mask = 16'hB8FF;
defparam \mem[117][67]~234 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[117][67]~235 (
	.dataa(\mem[117][67]~q ),
	.datab(\mem[117][67]~234_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[117]~q ),
	.cin(gnd),
	.combout(\mem[117][67]~235_combout ),
	.cout());
defparam \mem[117][67]~235 .lut_mask = 16'hEFFE;
defparam \mem[117][67]~235 .sum_lutc_input = "datac";

dffeas \mem[117][67] (
	.clk(clk),
	.d(\mem[117][67]~235_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[117][67]~q ),
	.prn(vcc));
defparam \mem[117][67] .is_wysiwyg = "true";
defparam \mem[117][67] .power_up = "low";

cycloneive_lcell_comb \mem[116][67]~232 (
	.dataa(\mem[117][67]~q ),
	.datab(\mem_used[117]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[116][67]~232_combout ),
	.cout());
defparam \mem[116][67]~232 .lut_mask = 16'hB8FF;
defparam \mem[116][67]~232 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[116][67]~233 (
	.dataa(\mem[116][67]~q ),
	.datab(\mem[116][67]~232_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[116]~q ),
	.cin(gnd),
	.combout(\mem[116][67]~233_combout ),
	.cout());
defparam \mem[116][67]~233 .lut_mask = 16'hEFFE;
defparam \mem[116][67]~233 .sum_lutc_input = "datac";

dffeas \mem[116][67] (
	.clk(clk),
	.d(\mem[116][67]~233_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[116][67]~q ),
	.prn(vcc));
defparam \mem[116][67] .is_wysiwyg = "true";
defparam \mem[116][67] .power_up = "low";

cycloneive_lcell_comb \mem[115][67]~230 (
	.dataa(\mem[116][67]~q ),
	.datab(\mem_used[116]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[115][67]~230_combout ),
	.cout());
defparam \mem[115][67]~230 .lut_mask = 16'hB8FF;
defparam \mem[115][67]~230 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[115][67]~231 (
	.dataa(\mem[115][67]~q ),
	.datab(\mem[115][67]~230_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[115]~q ),
	.cin(gnd),
	.combout(\mem[115][67]~231_combout ),
	.cout());
defparam \mem[115][67]~231 .lut_mask = 16'hEFFE;
defparam \mem[115][67]~231 .sum_lutc_input = "datac";

dffeas \mem[115][67] (
	.clk(clk),
	.d(\mem[115][67]~231_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[115][67]~q ),
	.prn(vcc));
defparam \mem[115][67] .is_wysiwyg = "true";
defparam \mem[115][67] .power_up = "low";

cycloneive_lcell_comb \mem[114][67]~228 (
	.dataa(\mem[115][67]~q ),
	.datab(\mem_used[115]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[114][67]~228_combout ),
	.cout());
defparam \mem[114][67]~228 .lut_mask = 16'hB8FF;
defparam \mem[114][67]~228 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[114][67]~229 (
	.dataa(\mem[114][67]~q ),
	.datab(\mem[114][67]~228_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[114]~q ),
	.cin(gnd),
	.combout(\mem[114][67]~229_combout ),
	.cout());
defparam \mem[114][67]~229 .lut_mask = 16'hEFFE;
defparam \mem[114][67]~229 .sum_lutc_input = "datac";

dffeas \mem[114][67] (
	.clk(clk),
	.d(\mem[114][67]~229_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[114][67]~q ),
	.prn(vcc));
defparam \mem[114][67] .is_wysiwyg = "true";
defparam \mem[114][67] .power_up = "low";

cycloneive_lcell_comb \mem[113][67]~226 (
	.dataa(\mem[114][67]~q ),
	.datab(\mem_used[114]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[113][67]~226_combout ),
	.cout());
defparam \mem[113][67]~226 .lut_mask = 16'hB8FF;
defparam \mem[113][67]~226 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[113][67]~227 (
	.dataa(\mem[113][67]~q ),
	.datab(\mem[113][67]~226_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[113]~q ),
	.cin(gnd),
	.combout(\mem[113][67]~227_combout ),
	.cout());
defparam \mem[113][67]~227 .lut_mask = 16'hEFFE;
defparam \mem[113][67]~227 .sum_lutc_input = "datac";

dffeas \mem[113][67] (
	.clk(clk),
	.d(\mem[113][67]~227_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[113][67]~q ),
	.prn(vcc));
defparam \mem[113][67] .is_wysiwyg = "true";
defparam \mem[113][67] .power_up = "low";

cycloneive_lcell_comb \mem[112][67]~224 (
	.dataa(\mem[113][67]~q ),
	.datab(\mem_used[113]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[112][67]~224_combout ),
	.cout());
defparam \mem[112][67]~224 .lut_mask = 16'hB8FF;
defparam \mem[112][67]~224 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[112][67]~225 (
	.dataa(\mem[112][67]~q ),
	.datab(\mem[112][67]~224_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[112]~q ),
	.cin(gnd),
	.combout(\mem[112][67]~225_combout ),
	.cout());
defparam \mem[112][67]~225 .lut_mask = 16'hEFFE;
defparam \mem[112][67]~225 .sum_lutc_input = "datac";

dffeas \mem[112][67] (
	.clk(clk),
	.d(\mem[112][67]~225_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[112][67]~q ),
	.prn(vcc));
defparam \mem[112][67] .is_wysiwyg = "true";
defparam \mem[112][67] .power_up = "low";

cycloneive_lcell_comb \mem[111][67]~222 (
	.dataa(\mem[112][67]~q ),
	.datab(\mem_used[112]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[111][67]~222_combout ),
	.cout());
defparam \mem[111][67]~222 .lut_mask = 16'hB8FF;
defparam \mem[111][67]~222 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[111][67]~223 (
	.dataa(\mem[111][67]~q ),
	.datab(\mem[111][67]~222_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[111]~q ),
	.cin(gnd),
	.combout(\mem[111][67]~223_combout ),
	.cout());
defparam \mem[111][67]~223 .lut_mask = 16'hEFFE;
defparam \mem[111][67]~223 .sum_lutc_input = "datac";

dffeas \mem[111][67] (
	.clk(clk),
	.d(\mem[111][67]~223_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[111][67]~q ),
	.prn(vcc));
defparam \mem[111][67] .is_wysiwyg = "true";
defparam \mem[111][67] .power_up = "low";

cycloneive_lcell_comb \mem[110][67]~220 (
	.dataa(\mem[111][67]~q ),
	.datab(\mem_used[111]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[110][67]~220_combout ),
	.cout());
defparam \mem[110][67]~220 .lut_mask = 16'hB8FF;
defparam \mem[110][67]~220 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[110][67]~221 (
	.dataa(\mem[110][67]~q ),
	.datab(\mem[110][67]~220_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[110]~q ),
	.cin(gnd),
	.combout(\mem[110][67]~221_combout ),
	.cout());
defparam \mem[110][67]~221 .lut_mask = 16'hEFFE;
defparam \mem[110][67]~221 .sum_lutc_input = "datac";

dffeas \mem[110][67] (
	.clk(clk),
	.d(\mem[110][67]~221_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[110][67]~q ),
	.prn(vcc));
defparam \mem[110][67] .is_wysiwyg = "true";
defparam \mem[110][67] .power_up = "low";

cycloneive_lcell_comb \mem[109][67]~218 (
	.dataa(\mem[110][67]~q ),
	.datab(\mem_used[110]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[109][67]~218_combout ),
	.cout());
defparam \mem[109][67]~218 .lut_mask = 16'hB8FF;
defparam \mem[109][67]~218 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[109][67]~219 (
	.dataa(\mem[109][67]~q ),
	.datab(\mem[109][67]~218_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[109]~q ),
	.cin(gnd),
	.combout(\mem[109][67]~219_combout ),
	.cout());
defparam \mem[109][67]~219 .lut_mask = 16'hEFFE;
defparam \mem[109][67]~219 .sum_lutc_input = "datac";

dffeas \mem[109][67] (
	.clk(clk),
	.d(\mem[109][67]~219_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[109][67]~q ),
	.prn(vcc));
defparam \mem[109][67] .is_wysiwyg = "true";
defparam \mem[109][67] .power_up = "low";

cycloneive_lcell_comb \mem[108][67]~216 (
	.dataa(\mem[109][67]~q ),
	.datab(\mem_used[109]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[108][67]~216_combout ),
	.cout());
defparam \mem[108][67]~216 .lut_mask = 16'hB8FF;
defparam \mem[108][67]~216 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[108][67]~217 (
	.dataa(\mem[108][67]~q ),
	.datab(\mem[108][67]~216_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[108]~q ),
	.cin(gnd),
	.combout(\mem[108][67]~217_combout ),
	.cout());
defparam \mem[108][67]~217 .lut_mask = 16'hEFFE;
defparam \mem[108][67]~217 .sum_lutc_input = "datac";

dffeas \mem[108][67] (
	.clk(clk),
	.d(\mem[108][67]~217_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[108][67]~q ),
	.prn(vcc));
defparam \mem[108][67] .is_wysiwyg = "true";
defparam \mem[108][67] .power_up = "low";

cycloneive_lcell_comb \mem[107][67]~214 (
	.dataa(\mem[108][67]~q ),
	.datab(\mem_used[108]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[107][67]~214_combout ),
	.cout());
defparam \mem[107][67]~214 .lut_mask = 16'hB8FF;
defparam \mem[107][67]~214 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[107][67]~215 (
	.dataa(\mem[107][67]~q ),
	.datab(\mem[107][67]~214_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[107]~q ),
	.cin(gnd),
	.combout(\mem[107][67]~215_combout ),
	.cout());
defparam \mem[107][67]~215 .lut_mask = 16'hEFFE;
defparam \mem[107][67]~215 .sum_lutc_input = "datac";

dffeas \mem[107][67] (
	.clk(clk),
	.d(\mem[107][67]~215_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[107][67]~q ),
	.prn(vcc));
defparam \mem[107][67] .is_wysiwyg = "true";
defparam \mem[107][67] .power_up = "low";

cycloneive_lcell_comb \mem[106][67]~212 (
	.dataa(\mem[107][67]~q ),
	.datab(\mem_used[107]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[106][67]~212_combout ),
	.cout());
defparam \mem[106][67]~212 .lut_mask = 16'hB8FF;
defparam \mem[106][67]~212 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[106][67]~213 (
	.dataa(\mem[106][67]~q ),
	.datab(\mem[106][67]~212_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[106]~q ),
	.cin(gnd),
	.combout(\mem[106][67]~213_combout ),
	.cout());
defparam \mem[106][67]~213 .lut_mask = 16'hEFFE;
defparam \mem[106][67]~213 .sum_lutc_input = "datac";

dffeas \mem[106][67] (
	.clk(clk),
	.d(\mem[106][67]~213_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[106][67]~q ),
	.prn(vcc));
defparam \mem[106][67] .is_wysiwyg = "true";
defparam \mem[106][67] .power_up = "low";

cycloneive_lcell_comb \mem[105][67]~210 (
	.dataa(\mem[106][67]~q ),
	.datab(\mem_used[106]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[105][67]~210_combout ),
	.cout());
defparam \mem[105][67]~210 .lut_mask = 16'hB8FF;
defparam \mem[105][67]~210 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[105][67]~211 (
	.dataa(\mem[105][67]~q ),
	.datab(\mem[105][67]~210_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[105]~q ),
	.cin(gnd),
	.combout(\mem[105][67]~211_combout ),
	.cout());
defparam \mem[105][67]~211 .lut_mask = 16'hEFFE;
defparam \mem[105][67]~211 .sum_lutc_input = "datac";

dffeas \mem[105][67] (
	.clk(clk),
	.d(\mem[105][67]~211_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[105][67]~q ),
	.prn(vcc));
defparam \mem[105][67] .is_wysiwyg = "true";
defparam \mem[105][67] .power_up = "low";

cycloneive_lcell_comb \mem[104][67]~208 (
	.dataa(\mem[105][67]~q ),
	.datab(\mem_used[105]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[104][67]~208_combout ),
	.cout());
defparam \mem[104][67]~208 .lut_mask = 16'hB8FF;
defparam \mem[104][67]~208 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[104][67]~209 (
	.dataa(\mem[104][67]~q ),
	.datab(\mem[104][67]~208_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[104]~q ),
	.cin(gnd),
	.combout(\mem[104][67]~209_combout ),
	.cout());
defparam \mem[104][67]~209 .lut_mask = 16'hEFFE;
defparam \mem[104][67]~209 .sum_lutc_input = "datac";

dffeas \mem[104][67] (
	.clk(clk),
	.d(\mem[104][67]~209_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[104][67]~q ),
	.prn(vcc));
defparam \mem[104][67] .is_wysiwyg = "true";
defparam \mem[104][67] .power_up = "low";

cycloneive_lcell_comb \mem[103][67]~206 (
	.dataa(\mem[104][67]~q ),
	.datab(\mem_used[104]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[103][67]~206_combout ),
	.cout());
defparam \mem[103][67]~206 .lut_mask = 16'hB8FF;
defparam \mem[103][67]~206 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[103][67]~207 (
	.dataa(\mem[103][67]~q ),
	.datab(\mem[103][67]~206_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[103]~q ),
	.cin(gnd),
	.combout(\mem[103][67]~207_combout ),
	.cout());
defparam \mem[103][67]~207 .lut_mask = 16'hEFFE;
defparam \mem[103][67]~207 .sum_lutc_input = "datac";

dffeas \mem[103][67] (
	.clk(clk),
	.d(\mem[103][67]~207_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[103][67]~q ),
	.prn(vcc));
defparam \mem[103][67] .is_wysiwyg = "true";
defparam \mem[103][67] .power_up = "low";

cycloneive_lcell_comb \mem[102][67]~204 (
	.dataa(\mem[103][67]~q ),
	.datab(\mem_used[103]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[102][67]~204_combout ),
	.cout());
defparam \mem[102][67]~204 .lut_mask = 16'hB8FF;
defparam \mem[102][67]~204 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[102][67]~205 (
	.dataa(\mem[102][67]~q ),
	.datab(\mem[102][67]~204_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[102]~q ),
	.cin(gnd),
	.combout(\mem[102][67]~205_combout ),
	.cout());
defparam \mem[102][67]~205 .lut_mask = 16'hEFFE;
defparam \mem[102][67]~205 .sum_lutc_input = "datac";

dffeas \mem[102][67] (
	.clk(clk),
	.d(\mem[102][67]~205_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[102][67]~q ),
	.prn(vcc));
defparam \mem[102][67] .is_wysiwyg = "true";
defparam \mem[102][67] .power_up = "low";

cycloneive_lcell_comb \mem[101][67]~202 (
	.dataa(\mem[102][67]~q ),
	.datab(\mem_used[102]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[101][67]~202_combout ),
	.cout());
defparam \mem[101][67]~202 .lut_mask = 16'hB8FF;
defparam \mem[101][67]~202 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[101][67]~203 (
	.dataa(\mem[101][67]~q ),
	.datab(\mem[101][67]~202_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[101]~q ),
	.cin(gnd),
	.combout(\mem[101][67]~203_combout ),
	.cout());
defparam \mem[101][67]~203 .lut_mask = 16'hEFFE;
defparam \mem[101][67]~203 .sum_lutc_input = "datac";

dffeas \mem[101][67] (
	.clk(clk),
	.d(\mem[101][67]~203_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[101][67]~q ),
	.prn(vcc));
defparam \mem[101][67] .is_wysiwyg = "true";
defparam \mem[101][67] .power_up = "low";

cycloneive_lcell_comb \mem[100][67]~200 (
	.dataa(\mem[101][67]~q ),
	.datab(\mem_used[101]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[100][67]~200_combout ),
	.cout());
defparam \mem[100][67]~200 .lut_mask = 16'hB8FF;
defparam \mem[100][67]~200 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[100][67]~201 (
	.dataa(\mem[100][67]~q ),
	.datab(\mem[100][67]~200_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[100]~q ),
	.cin(gnd),
	.combout(\mem[100][67]~201_combout ),
	.cout());
defparam \mem[100][67]~201 .lut_mask = 16'hEFFE;
defparam \mem[100][67]~201 .sum_lutc_input = "datac";

dffeas \mem[100][67] (
	.clk(clk),
	.d(\mem[100][67]~201_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[100][67]~q ),
	.prn(vcc));
defparam \mem[100][67] .is_wysiwyg = "true";
defparam \mem[100][67] .power_up = "low";

cycloneive_lcell_comb \mem[99][67]~198 (
	.dataa(\mem[100][67]~q ),
	.datab(\mem_used[100]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[99][67]~198_combout ),
	.cout());
defparam \mem[99][67]~198 .lut_mask = 16'hB8FF;
defparam \mem[99][67]~198 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[99][67]~199 (
	.dataa(\mem[99][67]~q ),
	.datab(\mem[99][67]~198_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[99]~q ),
	.cin(gnd),
	.combout(\mem[99][67]~199_combout ),
	.cout());
defparam \mem[99][67]~199 .lut_mask = 16'hEFFE;
defparam \mem[99][67]~199 .sum_lutc_input = "datac";

dffeas \mem[99][67] (
	.clk(clk),
	.d(\mem[99][67]~199_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[99][67]~q ),
	.prn(vcc));
defparam \mem[99][67] .is_wysiwyg = "true";
defparam \mem[99][67] .power_up = "low";

cycloneive_lcell_comb \mem[98][67]~196 (
	.dataa(\mem[99][67]~q ),
	.datab(\mem_used[99]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[98][67]~196_combout ),
	.cout());
defparam \mem[98][67]~196 .lut_mask = 16'hB8FF;
defparam \mem[98][67]~196 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[98][67]~197 (
	.dataa(\mem[98][67]~q ),
	.datab(\mem[98][67]~196_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[98]~q ),
	.cin(gnd),
	.combout(\mem[98][67]~197_combout ),
	.cout());
defparam \mem[98][67]~197 .lut_mask = 16'hEFFE;
defparam \mem[98][67]~197 .sum_lutc_input = "datac";

dffeas \mem[98][67] (
	.clk(clk),
	.d(\mem[98][67]~197_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[98][67]~q ),
	.prn(vcc));
defparam \mem[98][67] .is_wysiwyg = "true";
defparam \mem[98][67] .power_up = "low";

cycloneive_lcell_comb \mem[97][67]~194 (
	.dataa(\mem[98][67]~q ),
	.datab(\mem_used[98]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[97][67]~194_combout ),
	.cout());
defparam \mem[97][67]~194 .lut_mask = 16'hB8FF;
defparam \mem[97][67]~194 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[97][67]~195 (
	.dataa(\mem[97][67]~q ),
	.datab(\mem[97][67]~194_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[97]~q ),
	.cin(gnd),
	.combout(\mem[97][67]~195_combout ),
	.cout());
defparam \mem[97][67]~195 .lut_mask = 16'hEFFE;
defparam \mem[97][67]~195 .sum_lutc_input = "datac";

dffeas \mem[97][67] (
	.clk(clk),
	.d(\mem[97][67]~195_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[97][67]~q ),
	.prn(vcc));
defparam \mem[97][67] .is_wysiwyg = "true";
defparam \mem[97][67] .power_up = "low";

cycloneive_lcell_comb \mem[96][67]~192 (
	.dataa(\mem[97][67]~q ),
	.datab(\mem_used[97]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[96][67]~192_combout ),
	.cout());
defparam \mem[96][67]~192 .lut_mask = 16'hB8FF;
defparam \mem[96][67]~192 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[96][67]~193 (
	.dataa(\mem[96][67]~q ),
	.datab(\mem[96][67]~192_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[96]~q ),
	.cin(gnd),
	.combout(\mem[96][67]~193_combout ),
	.cout());
defparam \mem[96][67]~193 .lut_mask = 16'hEFFE;
defparam \mem[96][67]~193 .sum_lutc_input = "datac";

dffeas \mem[96][67] (
	.clk(clk),
	.d(\mem[96][67]~193_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[96][67]~q ),
	.prn(vcc));
defparam \mem[96][67] .is_wysiwyg = "true";
defparam \mem[96][67] .power_up = "low";

cycloneive_lcell_comb \mem[95][67]~190 (
	.dataa(\mem[96][67]~q ),
	.datab(\mem_used[96]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[95][67]~190_combout ),
	.cout());
defparam \mem[95][67]~190 .lut_mask = 16'hB8FF;
defparam \mem[95][67]~190 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[95][67]~191 (
	.dataa(\mem[95][67]~q ),
	.datab(\mem[95][67]~190_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[95]~q ),
	.cin(gnd),
	.combout(\mem[95][67]~191_combout ),
	.cout());
defparam \mem[95][67]~191 .lut_mask = 16'hEFFE;
defparam \mem[95][67]~191 .sum_lutc_input = "datac";

dffeas \mem[95][67] (
	.clk(clk),
	.d(\mem[95][67]~191_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[95][67]~q ),
	.prn(vcc));
defparam \mem[95][67] .is_wysiwyg = "true";
defparam \mem[95][67] .power_up = "low";

cycloneive_lcell_comb \mem[94][67]~188 (
	.dataa(\mem[95][67]~q ),
	.datab(\mem_used[95]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[94][67]~188_combout ),
	.cout());
defparam \mem[94][67]~188 .lut_mask = 16'hB8FF;
defparam \mem[94][67]~188 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[94][67]~189 (
	.dataa(\mem[94][67]~q ),
	.datab(\mem[94][67]~188_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[94]~q ),
	.cin(gnd),
	.combout(\mem[94][67]~189_combout ),
	.cout());
defparam \mem[94][67]~189 .lut_mask = 16'hEFFE;
defparam \mem[94][67]~189 .sum_lutc_input = "datac";

dffeas \mem[94][67] (
	.clk(clk),
	.d(\mem[94][67]~189_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[94][67]~q ),
	.prn(vcc));
defparam \mem[94][67] .is_wysiwyg = "true";
defparam \mem[94][67] .power_up = "low";

cycloneive_lcell_comb \mem[93][67]~186 (
	.dataa(\mem[94][67]~q ),
	.datab(\mem_used[94]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[93][67]~186_combout ),
	.cout());
defparam \mem[93][67]~186 .lut_mask = 16'hB8FF;
defparam \mem[93][67]~186 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[93][67]~187 (
	.dataa(\mem[93][67]~q ),
	.datab(\mem[93][67]~186_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[93]~q ),
	.cin(gnd),
	.combout(\mem[93][67]~187_combout ),
	.cout());
defparam \mem[93][67]~187 .lut_mask = 16'hEFFE;
defparam \mem[93][67]~187 .sum_lutc_input = "datac";

dffeas \mem[93][67] (
	.clk(clk),
	.d(\mem[93][67]~187_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[93][67]~q ),
	.prn(vcc));
defparam \mem[93][67] .is_wysiwyg = "true";
defparam \mem[93][67] .power_up = "low";

cycloneive_lcell_comb \mem[92][67]~184 (
	.dataa(\mem[93][67]~q ),
	.datab(\mem_used[93]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[92][67]~184_combout ),
	.cout());
defparam \mem[92][67]~184 .lut_mask = 16'hB8FF;
defparam \mem[92][67]~184 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[92][67]~185 (
	.dataa(\mem[92][67]~q ),
	.datab(\mem[92][67]~184_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[92]~q ),
	.cin(gnd),
	.combout(\mem[92][67]~185_combout ),
	.cout());
defparam \mem[92][67]~185 .lut_mask = 16'hEFFE;
defparam \mem[92][67]~185 .sum_lutc_input = "datac";

dffeas \mem[92][67] (
	.clk(clk),
	.d(\mem[92][67]~185_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[92][67]~q ),
	.prn(vcc));
defparam \mem[92][67] .is_wysiwyg = "true";
defparam \mem[92][67] .power_up = "low";

cycloneive_lcell_comb \mem[91][67]~182 (
	.dataa(\mem[92][67]~q ),
	.datab(\mem_used[92]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[91][67]~182_combout ),
	.cout());
defparam \mem[91][67]~182 .lut_mask = 16'hB8FF;
defparam \mem[91][67]~182 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[91][67]~183 (
	.dataa(\mem[91][67]~q ),
	.datab(\mem[91][67]~182_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[91]~q ),
	.cin(gnd),
	.combout(\mem[91][67]~183_combout ),
	.cout());
defparam \mem[91][67]~183 .lut_mask = 16'hEFFE;
defparam \mem[91][67]~183 .sum_lutc_input = "datac";

dffeas \mem[91][67] (
	.clk(clk),
	.d(\mem[91][67]~183_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[91][67]~q ),
	.prn(vcc));
defparam \mem[91][67] .is_wysiwyg = "true";
defparam \mem[91][67] .power_up = "low";

cycloneive_lcell_comb \mem[90][67]~180 (
	.dataa(\mem[91][67]~q ),
	.datab(\mem_used[91]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[90][67]~180_combout ),
	.cout());
defparam \mem[90][67]~180 .lut_mask = 16'hB8FF;
defparam \mem[90][67]~180 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[90][67]~181 (
	.dataa(\mem[90][67]~q ),
	.datab(\mem[90][67]~180_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[90]~q ),
	.cin(gnd),
	.combout(\mem[90][67]~181_combout ),
	.cout());
defparam \mem[90][67]~181 .lut_mask = 16'hEFFE;
defparam \mem[90][67]~181 .sum_lutc_input = "datac";

dffeas \mem[90][67] (
	.clk(clk),
	.d(\mem[90][67]~181_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[90][67]~q ),
	.prn(vcc));
defparam \mem[90][67] .is_wysiwyg = "true";
defparam \mem[90][67] .power_up = "low";

cycloneive_lcell_comb \mem[89][67]~178 (
	.dataa(\mem[90][67]~q ),
	.datab(\mem_used[90]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[89][67]~178_combout ),
	.cout());
defparam \mem[89][67]~178 .lut_mask = 16'hB8FF;
defparam \mem[89][67]~178 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[89][67]~179 (
	.dataa(\mem[89][67]~q ),
	.datab(\mem[89][67]~178_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[89]~q ),
	.cin(gnd),
	.combout(\mem[89][67]~179_combout ),
	.cout());
defparam \mem[89][67]~179 .lut_mask = 16'hEFFE;
defparam \mem[89][67]~179 .sum_lutc_input = "datac";

dffeas \mem[89][67] (
	.clk(clk),
	.d(\mem[89][67]~179_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[89][67]~q ),
	.prn(vcc));
defparam \mem[89][67] .is_wysiwyg = "true";
defparam \mem[89][67] .power_up = "low";

cycloneive_lcell_comb \mem[88][67]~176 (
	.dataa(\mem[89][67]~q ),
	.datab(\mem_used[89]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[88][67]~176_combout ),
	.cout());
defparam \mem[88][67]~176 .lut_mask = 16'hB8FF;
defparam \mem[88][67]~176 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[88][67]~177 (
	.dataa(\mem[88][67]~q ),
	.datab(\mem[88][67]~176_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[88]~q ),
	.cin(gnd),
	.combout(\mem[88][67]~177_combout ),
	.cout());
defparam \mem[88][67]~177 .lut_mask = 16'hEFFE;
defparam \mem[88][67]~177 .sum_lutc_input = "datac";

dffeas \mem[88][67] (
	.clk(clk),
	.d(\mem[88][67]~177_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[88][67]~q ),
	.prn(vcc));
defparam \mem[88][67] .is_wysiwyg = "true";
defparam \mem[88][67] .power_up = "low";

cycloneive_lcell_comb \mem[87][67]~174 (
	.dataa(\mem[88][67]~q ),
	.datab(\mem_used[88]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[87][67]~174_combout ),
	.cout());
defparam \mem[87][67]~174 .lut_mask = 16'hB8FF;
defparam \mem[87][67]~174 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[87][67]~175 (
	.dataa(\mem[87][67]~q ),
	.datab(\mem[87][67]~174_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[87]~q ),
	.cin(gnd),
	.combout(\mem[87][67]~175_combout ),
	.cout());
defparam \mem[87][67]~175 .lut_mask = 16'hEFFE;
defparam \mem[87][67]~175 .sum_lutc_input = "datac";

dffeas \mem[87][67] (
	.clk(clk),
	.d(\mem[87][67]~175_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[87][67]~q ),
	.prn(vcc));
defparam \mem[87][67] .is_wysiwyg = "true";
defparam \mem[87][67] .power_up = "low";

cycloneive_lcell_comb \mem[86][67]~172 (
	.dataa(\mem[87][67]~q ),
	.datab(\mem_used[87]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[86][67]~172_combout ),
	.cout());
defparam \mem[86][67]~172 .lut_mask = 16'hB8FF;
defparam \mem[86][67]~172 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[86][67]~173 (
	.dataa(\mem[86][67]~q ),
	.datab(\mem[86][67]~172_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[86]~q ),
	.cin(gnd),
	.combout(\mem[86][67]~173_combout ),
	.cout());
defparam \mem[86][67]~173 .lut_mask = 16'hEFFE;
defparam \mem[86][67]~173 .sum_lutc_input = "datac";

dffeas \mem[86][67] (
	.clk(clk),
	.d(\mem[86][67]~173_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[86][67]~q ),
	.prn(vcc));
defparam \mem[86][67] .is_wysiwyg = "true";
defparam \mem[86][67] .power_up = "low";

cycloneive_lcell_comb \mem[85][67]~170 (
	.dataa(\mem[86][67]~q ),
	.datab(\mem_used[86]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[85][67]~170_combout ),
	.cout());
defparam \mem[85][67]~170 .lut_mask = 16'hB8FF;
defparam \mem[85][67]~170 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[85][67]~171 (
	.dataa(\mem[85][67]~q ),
	.datab(\mem[85][67]~170_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[85]~q ),
	.cin(gnd),
	.combout(\mem[85][67]~171_combout ),
	.cout());
defparam \mem[85][67]~171 .lut_mask = 16'hEFFE;
defparam \mem[85][67]~171 .sum_lutc_input = "datac";

dffeas \mem[85][67] (
	.clk(clk),
	.d(\mem[85][67]~171_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[85][67]~q ),
	.prn(vcc));
defparam \mem[85][67] .is_wysiwyg = "true";
defparam \mem[85][67] .power_up = "low";

cycloneive_lcell_comb \mem[84][67]~168 (
	.dataa(\mem[85][67]~q ),
	.datab(\mem_used[85]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[84][67]~168_combout ),
	.cout());
defparam \mem[84][67]~168 .lut_mask = 16'hB8FF;
defparam \mem[84][67]~168 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[84][67]~169 (
	.dataa(\mem[84][67]~q ),
	.datab(\mem[84][67]~168_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[84]~q ),
	.cin(gnd),
	.combout(\mem[84][67]~169_combout ),
	.cout());
defparam \mem[84][67]~169 .lut_mask = 16'hEFFE;
defparam \mem[84][67]~169 .sum_lutc_input = "datac";

dffeas \mem[84][67] (
	.clk(clk),
	.d(\mem[84][67]~169_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[84][67]~q ),
	.prn(vcc));
defparam \mem[84][67] .is_wysiwyg = "true";
defparam \mem[84][67] .power_up = "low";

cycloneive_lcell_comb \mem[83][67]~166 (
	.dataa(\mem[84][67]~q ),
	.datab(\mem_used[84]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[83][67]~166_combout ),
	.cout());
defparam \mem[83][67]~166 .lut_mask = 16'hB8FF;
defparam \mem[83][67]~166 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[83][67]~167 (
	.dataa(\mem[83][67]~q ),
	.datab(\mem[83][67]~166_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[83]~q ),
	.cin(gnd),
	.combout(\mem[83][67]~167_combout ),
	.cout());
defparam \mem[83][67]~167 .lut_mask = 16'hEFFE;
defparam \mem[83][67]~167 .sum_lutc_input = "datac";

dffeas \mem[83][67] (
	.clk(clk),
	.d(\mem[83][67]~167_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[83][67]~q ),
	.prn(vcc));
defparam \mem[83][67] .is_wysiwyg = "true";
defparam \mem[83][67] .power_up = "low";

cycloneive_lcell_comb \mem[82][67]~164 (
	.dataa(\mem[83][67]~q ),
	.datab(\mem_used[83]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[82][67]~164_combout ),
	.cout());
defparam \mem[82][67]~164 .lut_mask = 16'hB8FF;
defparam \mem[82][67]~164 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[82][67]~165 (
	.dataa(\mem[82][67]~q ),
	.datab(\mem[82][67]~164_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[82]~q ),
	.cin(gnd),
	.combout(\mem[82][67]~165_combout ),
	.cout());
defparam \mem[82][67]~165 .lut_mask = 16'hEFFE;
defparam \mem[82][67]~165 .sum_lutc_input = "datac";

dffeas \mem[82][67] (
	.clk(clk),
	.d(\mem[82][67]~165_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[82][67]~q ),
	.prn(vcc));
defparam \mem[82][67] .is_wysiwyg = "true";
defparam \mem[82][67] .power_up = "low";

cycloneive_lcell_comb \mem[81][67]~162 (
	.dataa(\mem[82][67]~q ),
	.datab(\mem_used[82]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[81][67]~162_combout ),
	.cout());
defparam \mem[81][67]~162 .lut_mask = 16'hB8FF;
defparam \mem[81][67]~162 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[81][67]~163 (
	.dataa(\mem[81][67]~q ),
	.datab(\mem[81][67]~162_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[81]~q ),
	.cin(gnd),
	.combout(\mem[81][67]~163_combout ),
	.cout());
defparam \mem[81][67]~163 .lut_mask = 16'hEFFE;
defparam \mem[81][67]~163 .sum_lutc_input = "datac";

dffeas \mem[81][67] (
	.clk(clk),
	.d(\mem[81][67]~163_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[81][67]~q ),
	.prn(vcc));
defparam \mem[81][67] .is_wysiwyg = "true";
defparam \mem[81][67] .power_up = "low";

cycloneive_lcell_comb \mem[80][67]~160 (
	.dataa(\mem[81][67]~q ),
	.datab(\mem_used[81]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[80][67]~160_combout ),
	.cout());
defparam \mem[80][67]~160 .lut_mask = 16'hB8FF;
defparam \mem[80][67]~160 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[80][67]~161 (
	.dataa(\mem[80][67]~q ),
	.datab(\mem[80][67]~160_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[80]~q ),
	.cin(gnd),
	.combout(\mem[80][67]~161_combout ),
	.cout());
defparam \mem[80][67]~161 .lut_mask = 16'hEFFE;
defparam \mem[80][67]~161 .sum_lutc_input = "datac";

dffeas \mem[80][67] (
	.clk(clk),
	.d(\mem[80][67]~161_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[80][67]~q ),
	.prn(vcc));
defparam \mem[80][67] .is_wysiwyg = "true";
defparam \mem[80][67] .power_up = "low";

cycloneive_lcell_comb \mem[79][67]~158 (
	.dataa(\mem[80][67]~q ),
	.datab(\mem_used[80]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[79][67]~158_combout ),
	.cout());
defparam \mem[79][67]~158 .lut_mask = 16'hB8FF;
defparam \mem[79][67]~158 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[79][67]~159 (
	.dataa(\mem[79][67]~q ),
	.datab(\mem[79][67]~158_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[79]~q ),
	.cin(gnd),
	.combout(\mem[79][67]~159_combout ),
	.cout());
defparam \mem[79][67]~159 .lut_mask = 16'hEFFE;
defparam \mem[79][67]~159 .sum_lutc_input = "datac";

dffeas \mem[79][67] (
	.clk(clk),
	.d(\mem[79][67]~159_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[79][67]~q ),
	.prn(vcc));
defparam \mem[79][67] .is_wysiwyg = "true";
defparam \mem[79][67] .power_up = "low";

cycloneive_lcell_comb \mem[78][67]~156 (
	.dataa(\mem[79][67]~q ),
	.datab(\mem_used[79]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[78][67]~156_combout ),
	.cout());
defparam \mem[78][67]~156 .lut_mask = 16'hB8FF;
defparam \mem[78][67]~156 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[78][67]~157 (
	.dataa(\mem[78][67]~q ),
	.datab(\mem[78][67]~156_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[78]~q ),
	.cin(gnd),
	.combout(\mem[78][67]~157_combout ),
	.cout());
defparam \mem[78][67]~157 .lut_mask = 16'hEFFE;
defparam \mem[78][67]~157 .sum_lutc_input = "datac";

dffeas \mem[78][67] (
	.clk(clk),
	.d(\mem[78][67]~157_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[78][67]~q ),
	.prn(vcc));
defparam \mem[78][67] .is_wysiwyg = "true";
defparam \mem[78][67] .power_up = "low";

cycloneive_lcell_comb \mem[77][67]~154 (
	.dataa(\mem[78][67]~q ),
	.datab(\mem_used[78]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[77][67]~154_combout ),
	.cout());
defparam \mem[77][67]~154 .lut_mask = 16'hB8FF;
defparam \mem[77][67]~154 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[77][67]~155 (
	.dataa(\mem[77][67]~q ),
	.datab(\mem[77][67]~154_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[77]~q ),
	.cin(gnd),
	.combout(\mem[77][67]~155_combout ),
	.cout());
defparam \mem[77][67]~155 .lut_mask = 16'hEFFE;
defparam \mem[77][67]~155 .sum_lutc_input = "datac";

dffeas \mem[77][67] (
	.clk(clk),
	.d(\mem[77][67]~155_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[77][67]~q ),
	.prn(vcc));
defparam \mem[77][67] .is_wysiwyg = "true";
defparam \mem[77][67] .power_up = "low";

cycloneive_lcell_comb \mem[76][67]~152 (
	.dataa(\mem[77][67]~q ),
	.datab(\mem_used[77]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[76][67]~152_combout ),
	.cout());
defparam \mem[76][67]~152 .lut_mask = 16'hB8FF;
defparam \mem[76][67]~152 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[76][67]~153 (
	.dataa(\mem[76][67]~q ),
	.datab(\mem[76][67]~152_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[76]~q ),
	.cin(gnd),
	.combout(\mem[76][67]~153_combout ),
	.cout());
defparam \mem[76][67]~153 .lut_mask = 16'hEFFE;
defparam \mem[76][67]~153 .sum_lutc_input = "datac";

dffeas \mem[76][67] (
	.clk(clk),
	.d(\mem[76][67]~153_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[76][67]~q ),
	.prn(vcc));
defparam \mem[76][67] .is_wysiwyg = "true";
defparam \mem[76][67] .power_up = "low";

cycloneive_lcell_comb \mem[75][67]~150 (
	.dataa(\mem[76][67]~q ),
	.datab(\mem_used[76]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[75][67]~150_combout ),
	.cout());
defparam \mem[75][67]~150 .lut_mask = 16'hB8FF;
defparam \mem[75][67]~150 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[75][67]~151 (
	.dataa(\mem[75][67]~q ),
	.datab(\mem[75][67]~150_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[75]~q ),
	.cin(gnd),
	.combout(\mem[75][67]~151_combout ),
	.cout());
defparam \mem[75][67]~151 .lut_mask = 16'hEFFE;
defparam \mem[75][67]~151 .sum_lutc_input = "datac";

dffeas \mem[75][67] (
	.clk(clk),
	.d(\mem[75][67]~151_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[75][67]~q ),
	.prn(vcc));
defparam \mem[75][67] .is_wysiwyg = "true";
defparam \mem[75][67] .power_up = "low";

cycloneive_lcell_comb \mem[74][67]~148 (
	.dataa(\mem[75][67]~q ),
	.datab(\mem_used[75]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[74][67]~148_combout ),
	.cout());
defparam \mem[74][67]~148 .lut_mask = 16'hB8FF;
defparam \mem[74][67]~148 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[74][67]~149 (
	.dataa(\mem[74][67]~q ),
	.datab(\mem[74][67]~148_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[74]~q ),
	.cin(gnd),
	.combout(\mem[74][67]~149_combout ),
	.cout());
defparam \mem[74][67]~149 .lut_mask = 16'hEFFE;
defparam \mem[74][67]~149 .sum_lutc_input = "datac";

dffeas \mem[74][67] (
	.clk(clk),
	.d(\mem[74][67]~149_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[74][67]~q ),
	.prn(vcc));
defparam \mem[74][67] .is_wysiwyg = "true";
defparam \mem[74][67] .power_up = "low";

cycloneive_lcell_comb \mem[73][67]~146 (
	.dataa(\mem[74][67]~q ),
	.datab(\mem_used[74]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[73][67]~146_combout ),
	.cout());
defparam \mem[73][67]~146 .lut_mask = 16'hB8FF;
defparam \mem[73][67]~146 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[73][67]~147 (
	.dataa(\mem[73][67]~q ),
	.datab(\mem[73][67]~146_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[73]~q ),
	.cin(gnd),
	.combout(\mem[73][67]~147_combout ),
	.cout());
defparam \mem[73][67]~147 .lut_mask = 16'hEFFE;
defparam \mem[73][67]~147 .sum_lutc_input = "datac";

dffeas \mem[73][67] (
	.clk(clk),
	.d(\mem[73][67]~147_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[73][67]~q ),
	.prn(vcc));
defparam \mem[73][67] .is_wysiwyg = "true";
defparam \mem[73][67] .power_up = "low";

cycloneive_lcell_comb \mem[72][67]~144 (
	.dataa(\mem[73][67]~q ),
	.datab(\mem_used[73]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[72][67]~144_combout ),
	.cout());
defparam \mem[72][67]~144 .lut_mask = 16'hB8FF;
defparam \mem[72][67]~144 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[72][67]~145 (
	.dataa(\mem[72][67]~q ),
	.datab(\mem[72][67]~144_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[72]~q ),
	.cin(gnd),
	.combout(\mem[72][67]~145_combout ),
	.cout());
defparam \mem[72][67]~145 .lut_mask = 16'hEFFE;
defparam \mem[72][67]~145 .sum_lutc_input = "datac";

dffeas \mem[72][67] (
	.clk(clk),
	.d(\mem[72][67]~145_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[72][67]~q ),
	.prn(vcc));
defparam \mem[72][67] .is_wysiwyg = "true";
defparam \mem[72][67] .power_up = "low";

cycloneive_lcell_comb \mem[71][67]~142 (
	.dataa(\mem[72][67]~q ),
	.datab(\mem_used[72]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[71][67]~142_combout ),
	.cout());
defparam \mem[71][67]~142 .lut_mask = 16'hB8FF;
defparam \mem[71][67]~142 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[71][67]~143 (
	.dataa(\mem[71][67]~q ),
	.datab(\mem[71][67]~142_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[71]~q ),
	.cin(gnd),
	.combout(\mem[71][67]~143_combout ),
	.cout());
defparam \mem[71][67]~143 .lut_mask = 16'hEFFE;
defparam \mem[71][67]~143 .sum_lutc_input = "datac";

dffeas \mem[71][67] (
	.clk(clk),
	.d(\mem[71][67]~143_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[71][67]~q ),
	.prn(vcc));
defparam \mem[71][67] .is_wysiwyg = "true";
defparam \mem[71][67] .power_up = "low";

cycloneive_lcell_comb \mem[70][67]~140 (
	.dataa(\mem[71][67]~q ),
	.datab(\mem_used[71]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[70][67]~140_combout ),
	.cout());
defparam \mem[70][67]~140 .lut_mask = 16'hB8FF;
defparam \mem[70][67]~140 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[70][67]~141 (
	.dataa(\mem[70][67]~q ),
	.datab(\mem[70][67]~140_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[70]~q ),
	.cin(gnd),
	.combout(\mem[70][67]~141_combout ),
	.cout());
defparam \mem[70][67]~141 .lut_mask = 16'hEFFE;
defparam \mem[70][67]~141 .sum_lutc_input = "datac";

dffeas \mem[70][67] (
	.clk(clk),
	.d(\mem[70][67]~141_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[70][67]~q ),
	.prn(vcc));
defparam \mem[70][67] .is_wysiwyg = "true";
defparam \mem[70][67] .power_up = "low";

cycloneive_lcell_comb \mem[69][67]~138 (
	.dataa(\mem[70][67]~q ),
	.datab(\mem_used[70]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[69][67]~138_combout ),
	.cout());
defparam \mem[69][67]~138 .lut_mask = 16'hB8FF;
defparam \mem[69][67]~138 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[69][67]~139 (
	.dataa(\mem[69][67]~q ),
	.datab(\mem[69][67]~138_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[69]~q ),
	.cin(gnd),
	.combout(\mem[69][67]~139_combout ),
	.cout());
defparam \mem[69][67]~139 .lut_mask = 16'hEFFE;
defparam \mem[69][67]~139 .sum_lutc_input = "datac";

dffeas \mem[69][67] (
	.clk(clk),
	.d(\mem[69][67]~139_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[69][67]~q ),
	.prn(vcc));
defparam \mem[69][67] .is_wysiwyg = "true";
defparam \mem[69][67] .power_up = "low";

cycloneive_lcell_comb \mem[68][67]~136 (
	.dataa(\mem[69][67]~q ),
	.datab(\mem_used[69]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[68][67]~136_combout ),
	.cout());
defparam \mem[68][67]~136 .lut_mask = 16'hB8FF;
defparam \mem[68][67]~136 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[68][67]~137 (
	.dataa(\mem[68][67]~q ),
	.datab(\mem[68][67]~136_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[68]~q ),
	.cin(gnd),
	.combout(\mem[68][67]~137_combout ),
	.cout());
defparam \mem[68][67]~137 .lut_mask = 16'hEFFE;
defparam \mem[68][67]~137 .sum_lutc_input = "datac";

dffeas \mem[68][67] (
	.clk(clk),
	.d(\mem[68][67]~137_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[68][67]~q ),
	.prn(vcc));
defparam \mem[68][67] .is_wysiwyg = "true";
defparam \mem[68][67] .power_up = "low";

cycloneive_lcell_comb \mem[67][67]~134 (
	.dataa(\mem[68][67]~q ),
	.datab(\mem_used[68]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[67][67]~134_combout ),
	.cout());
defparam \mem[67][67]~134 .lut_mask = 16'hB8FF;
defparam \mem[67][67]~134 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[67][67]~135 (
	.dataa(\mem[67][67]~q ),
	.datab(\mem[67][67]~134_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[67]~q ),
	.cin(gnd),
	.combout(\mem[67][67]~135_combout ),
	.cout());
defparam \mem[67][67]~135 .lut_mask = 16'hEFFE;
defparam \mem[67][67]~135 .sum_lutc_input = "datac";

dffeas \mem[67][67] (
	.clk(clk),
	.d(\mem[67][67]~135_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[67][67]~q ),
	.prn(vcc));
defparam \mem[67][67] .is_wysiwyg = "true";
defparam \mem[67][67] .power_up = "low";

cycloneive_lcell_comb \mem[66][67]~132 (
	.dataa(\mem[67][67]~q ),
	.datab(\mem_used[67]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[66][67]~132_combout ),
	.cout());
defparam \mem[66][67]~132 .lut_mask = 16'hB8FF;
defparam \mem[66][67]~132 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[66][67]~133 (
	.dataa(\mem[66][67]~q ),
	.datab(\mem[66][67]~132_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[66]~q ),
	.cin(gnd),
	.combout(\mem[66][67]~133_combout ),
	.cout());
defparam \mem[66][67]~133 .lut_mask = 16'hEFFE;
defparam \mem[66][67]~133 .sum_lutc_input = "datac";

dffeas \mem[66][67] (
	.clk(clk),
	.d(\mem[66][67]~133_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[66][67]~q ),
	.prn(vcc));
defparam \mem[66][67] .is_wysiwyg = "true";
defparam \mem[66][67] .power_up = "low";

cycloneive_lcell_comb \mem[65][67]~130 (
	.dataa(\mem[66][67]~q ),
	.datab(\mem_used[66]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[65][67]~130_combout ),
	.cout());
defparam \mem[65][67]~130 .lut_mask = 16'hB8FF;
defparam \mem[65][67]~130 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[65][67]~131 (
	.dataa(\mem[65][67]~q ),
	.datab(\mem[65][67]~130_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[65]~q ),
	.cin(gnd),
	.combout(\mem[65][67]~131_combout ),
	.cout());
defparam \mem[65][67]~131 .lut_mask = 16'hEFFE;
defparam \mem[65][67]~131 .sum_lutc_input = "datac";

dffeas \mem[65][67] (
	.clk(clk),
	.d(\mem[65][67]~131_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[65][67]~q ),
	.prn(vcc));
defparam \mem[65][67] .is_wysiwyg = "true";
defparam \mem[65][67] .power_up = "low";

cycloneive_lcell_comb \mem[64][67]~128 (
	.dataa(\mem[65][67]~q ),
	.datab(\mem_used[65]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[64][67]~128_combout ),
	.cout());
defparam \mem[64][67]~128 .lut_mask = 16'hB8FF;
defparam \mem[64][67]~128 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[64][67]~129 (
	.dataa(\mem[64][67]~q ),
	.datab(\mem[64][67]~128_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[64]~q ),
	.cin(gnd),
	.combout(\mem[64][67]~129_combout ),
	.cout());
defparam \mem[64][67]~129 .lut_mask = 16'hEFFE;
defparam \mem[64][67]~129 .sum_lutc_input = "datac";

dffeas \mem[64][67] (
	.clk(clk),
	.d(\mem[64][67]~129_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[64][67]~q ),
	.prn(vcc));
defparam \mem[64][67] .is_wysiwyg = "true";
defparam \mem[64][67] .power_up = "low";

cycloneive_lcell_comb \mem[63][67]~126 (
	.dataa(\mem[64][67]~q ),
	.datab(\mem_used[64]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[63][67]~126_combout ),
	.cout());
defparam \mem[63][67]~126 .lut_mask = 16'hB8FF;
defparam \mem[63][67]~126 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[63][67]~127 (
	.dataa(\mem[63][67]~q ),
	.datab(\mem[63][67]~126_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[63]~q ),
	.cin(gnd),
	.combout(\mem[63][67]~127_combout ),
	.cout());
defparam \mem[63][67]~127 .lut_mask = 16'hEFFE;
defparam \mem[63][67]~127 .sum_lutc_input = "datac";

dffeas \mem[63][67] (
	.clk(clk),
	.d(\mem[63][67]~127_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[63][67]~q ),
	.prn(vcc));
defparam \mem[63][67] .is_wysiwyg = "true";
defparam \mem[63][67] .power_up = "low";

cycloneive_lcell_comb \mem[62][67]~124 (
	.dataa(\mem[63][67]~q ),
	.datab(\mem_used[63]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[62][67]~124_combout ),
	.cout());
defparam \mem[62][67]~124 .lut_mask = 16'hB8FF;
defparam \mem[62][67]~124 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[62][67]~125 (
	.dataa(\mem[62][67]~q ),
	.datab(\mem[62][67]~124_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[62]~q ),
	.cin(gnd),
	.combout(\mem[62][67]~125_combout ),
	.cout());
defparam \mem[62][67]~125 .lut_mask = 16'hEFFE;
defparam \mem[62][67]~125 .sum_lutc_input = "datac";

dffeas \mem[62][67] (
	.clk(clk),
	.d(\mem[62][67]~125_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[62][67]~q ),
	.prn(vcc));
defparam \mem[62][67] .is_wysiwyg = "true";
defparam \mem[62][67] .power_up = "low";

cycloneive_lcell_comb \mem[61][67]~122 (
	.dataa(\mem[62][67]~q ),
	.datab(\mem_used[62]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[61][67]~122_combout ),
	.cout());
defparam \mem[61][67]~122 .lut_mask = 16'hB8FF;
defparam \mem[61][67]~122 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[61][67]~123 (
	.dataa(\mem[61][67]~q ),
	.datab(\mem[61][67]~122_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[61]~q ),
	.cin(gnd),
	.combout(\mem[61][67]~123_combout ),
	.cout());
defparam \mem[61][67]~123 .lut_mask = 16'hEFFE;
defparam \mem[61][67]~123 .sum_lutc_input = "datac";

dffeas \mem[61][67] (
	.clk(clk),
	.d(\mem[61][67]~123_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[61][67]~q ),
	.prn(vcc));
defparam \mem[61][67] .is_wysiwyg = "true";
defparam \mem[61][67] .power_up = "low";

cycloneive_lcell_comb \mem[60][67]~120 (
	.dataa(\mem[61][67]~q ),
	.datab(\mem_used[61]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[60][67]~120_combout ),
	.cout());
defparam \mem[60][67]~120 .lut_mask = 16'hB8FF;
defparam \mem[60][67]~120 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[60][67]~121 (
	.dataa(\mem[60][67]~q ),
	.datab(\mem[60][67]~120_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[60]~q ),
	.cin(gnd),
	.combout(\mem[60][67]~121_combout ),
	.cout());
defparam \mem[60][67]~121 .lut_mask = 16'hEFFE;
defparam \mem[60][67]~121 .sum_lutc_input = "datac";

dffeas \mem[60][67] (
	.clk(clk),
	.d(\mem[60][67]~121_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[60][67]~q ),
	.prn(vcc));
defparam \mem[60][67] .is_wysiwyg = "true";
defparam \mem[60][67] .power_up = "low";

cycloneive_lcell_comb \mem[59][67]~118 (
	.dataa(\mem[60][67]~q ),
	.datab(\mem_used[60]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[59][67]~118_combout ),
	.cout());
defparam \mem[59][67]~118 .lut_mask = 16'hB8FF;
defparam \mem[59][67]~118 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[59][67]~119 (
	.dataa(\mem[59][67]~q ),
	.datab(\mem[59][67]~118_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[59]~q ),
	.cin(gnd),
	.combout(\mem[59][67]~119_combout ),
	.cout());
defparam \mem[59][67]~119 .lut_mask = 16'hEFFE;
defparam \mem[59][67]~119 .sum_lutc_input = "datac";

dffeas \mem[59][67] (
	.clk(clk),
	.d(\mem[59][67]~119_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[59][67]~q ),
	.prn(vcc));
defparam \mem[59][67] .is_wysiwyg = "true";
defparam \mem[59][67] .power_up = "low";

cycloneive_lcell_comb \mem[58][67]~116 (
	.dataa(\mem[59][67]~q ),
	.datab(\mem_used[59]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[58][67]~116_combout ),
	.cout());
defparam \mem[58][67]~116 .lut_mask = 16'hB8FF;
defparam \mem[58][67]~116 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[58][67]~117 (
	.dataa(\mem[58][67]~q ),
	.datab(\mem[58][67]~116_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[58]~q ),
	.cin(gnd),
	.combout(\mem[58][67]~117_combout ),
	.cout());
defparam \mem[58][67]~117 .lut_mask = 16'hEFFE;
defparam \mem[58][67]~117 .sum_lutc_input = "datac";

dffeas \mem[58][67] (
	.clk(clk),
	.d(\mem[58][67]~117_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[58][67]~q ),
	.prn(vcc));
defparam \mem[58][67] .is_wysiwyg = "true";
defparam \mem[58][67] .power_up = "low";

cycloneive_lcell_comb \mem[57][67]~114 (
	.dataa(\mem[58][67]~q ),
	.datab(\mem_used[58]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[57][67]~114_combout ),
	.cout());
defparam \mem[57][67]~114 .lut_mask = 16'hB8FF;
defparam \mem[57][67]~114 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[57][67]~115 (
	.dataa(\mem[57][67]~q ),
	.datab(\mem[57][67]~114_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[57]~q ),
	.cin(gnd),
	.combout(\mem[57][67]~115_combout ),
	.cout());
defparam \mem[57][67]~115 .lut_mask = 16'hEFFE;
defparam \mem[57][67]~115 .sum_lutc_input = "datac";

dffeas \mem[57][67] (
	.clk(clk),
	.d(\mem[57][67]~115_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[57][67]~q ),
	.prn(vcc));
defparam \mem[57][67] .is_wysiwyg = "true";
defparam \mem[57][67] .power_up = "low";

cycloneive_lcell_comb \mem[56][67]~112 (
	.dataa(\mem[57][67]~q ),
	.datab(\mem_used[57]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[56][67]~112_combout ),
	.cout());
defparam \mem[56][67]~112 .lut_mask = 16'hB8FF;
defparam \mem[56][67]~112 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[56][67]~113 (
	.dataa(\mem[56][67]~q ),
	.datab(\mem[56][67]~112_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[56]~q ),
	.cin(gnd),
	.combout(\mem[56][67]~113_combout ),
	.cout());
defparam \mem[56][67]~113 .lut_mask = 16'hEFFE;
defparam \mem[56][67]~113 .sum_lutc_input = "datac";

dffeas \mem[56][67] (
	.clk(clk),
	.d(\mem[56][67]~113_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[56][67]~q ),
	.prn(vcc));
defparam \mem[56][67] .is_wysiwyg = "true";
defparam \mem[56][67] .power_up = "low";

cycloneive_lcell_comb \mem[55][67]~110 (
	.dataa(\mem[56][67]~q ),
	.datab(\mem_used[56]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[55][67]~110_combout ),
	.cout());
defparam \mem[55][67]~110 .lut_mask = 16'hB8FF;
defparam \mem[55][67]~110 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[55][67]~111 (
	.dataa(\mem[55][67]~q ),
	.datab(\mem[55][67]~110_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[55]~q ),
	.cin(gnd),
	.combout(\mem[55][67]~111_combout ),
	.cout());
defparam \mem[55][67]~111 .lut_mask = 16'hEFFE;
defparam \mem[55][67]~111 .sum_lutc_input = "datac";

dffeas \mem[55][67] (
	.clk(clk),
	.d(\mem[55][67]~111_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[55][67]~q ),
	.prn(vcc));
defparam \mem[55][67] .is_wysiwyg = "true";
defparam \mem[55][67] .power_up = "low";

cycloneive_lcell_comb \mem[54][67]~108 (
	.dataa(\mem[55][67]~q ),
	.datab(\mem_used[55]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[54][67]~108_combout ),
	.cout());
defparam \mem[54][67]~108 .lut_mask = 16'hB8FF;
defparam \mem[54][67]~108 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[54][67]~109 (
	.dataa(\mem[54][67]~q ),
	.datab(\mem[54][67]~108_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[54]~q ),
	.cin(gnd),
	.combout(\mem[54][67]~109_combout ),
	.cout());
defparam \mem[54][67]~109 .lut_mask = 16'hEFFE;
defparam \mem[54][67]~109 .sum_lutc_input = "datac";

dffeas \mem[54][67] (
	.clk(clk),
	.d(\mem[54][67]~109_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[54][67]~q ),
	.prn(vcc));
defparam \mem[54][67] .is_wysiwyg = "true";
defparam \mem[54][67] .power_up = "low";

cycloneive_lcell_comb \mem[53][67]~106 (
	.dataa(\mem[54][67]~q ),
	.datab(\mem_used[54]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[53][67]~106_combout ),
	.cout());
defparam \mem[53][67]~106 .lut_mask = 16'hB8FF;
defparam \mem[53][67]~106 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[53][67]~107 (
	.dataa(\mem[53][67]~q ),
	.datab(\mem[53][67]~106_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[53]~q ),
	.cin(gnd),
	.combout(\mem[53][67]~107_combout ),
	.cout());
defparam \mem[53][67]~107 .lut_mask = 16'hEFFE;
defparam \mem[53][67]~107 .sum_lutc_input = "datac";

dffeas \mem[53][67] (
	.clk(clk),
	.d(\mem[53][67]~107_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[53][67]~q ),
	.prn(vcc));
defparam \mem[53][67] .is_wysiwyg = "true";
defparam \mem[53][67] .power_up = "low";

cycloneive_lcell_comb \mem[52][67]~104 (
	.dataa(\mem[53][67]~q ),
	.datab(\mem_used[53]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[52][67]~104_combout ),
	.cout());
defparam \mem[52][67]~104 .lut_mask = 16'hB8FF;
defparam \mem[52][67]~104 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[52][67]~105 (
	.dataa(\mem[52][67]~q ),
	.datab(\mem[52][67]~104_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[52]~q ),
	.cin(gnd),
	.combout(\mem[52][67]~105_combout ),
	.cout());
defparam \mem[52][67]~105 .lut_mask = 16'hEFFE;
defparam \mem[52][67]~105 .sum_lutc_input = "datac";

dffeas \mem[52][67] (
	.clk(clk),
	.d(\mem[52][67]~105_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[52][67]~q ),
	.prn(vcc));
defparam \mem[52][67] .is_wysiwyg = "true";
defparam \mem[52][67] .power_up = "low";

cycloneive_lcell_comb \mem[51][67]~102 (
	.dataa(\mem[52][67]~q ),
	.datab(\mem_used[52]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[51][67]~102_combout ),
	.cout());
defparam \mem[51][67]~102 .lut_mask = 16'hB8FF;
defparam \mem[51][67]~102 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[51][67]~103 (
	.dataa(\mem[51][67]~q ),
	.datab(\mem[51][67]~102_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[51]~q ),
	.cin(gnd),
	.combout(\mem[51][67]~103_combout ),
	.cout());
defparam \mem[51][67]~103 .lut_mask = 16'hEFFE;
defparam \mem[51][67]~103 .sum_lutc_input = "datac";

dffeas \mem[51][67] (
	.clk(clk),
	.d(\mem[51][67]~103_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[51][67]~q ),
	.prn(vcc));
defparam \mem[51][67] .is_wysiwyg = "true";
defparam \mem[51][67] .power_up = "low";

cycloneive_lcell_comb \mem[50][67]~100 (
	.dataa(\mem[51][67]~q ),
	.datab(\mem_used[51]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[50][67]~100_combout ),
	.cout());
defparam \mem[50][67]~100 .lut_mask = 16'hB8FF;
defparam \mem[50][67]~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[50][67]~101 (
	.dataa(\mem[50][67]~q ),
	.datab(\mem[50][67]~100_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[50]~q ),
	.cin(gnd),
	.combout(\mem[50][67]~101_combout ),
	.cout());
defparam \mem[50][67]~101 .lut_mask = 16'hEFFE;
defparam \mem[50][67]~101 .sum_lutc_input = "datac";

dffeas \mem[50][67] (
	.clk(clk),
	.d(\mem[50][67]~101_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[50][67]~q ),
	.prn(vcc));
defparam \mem[50][67] .is_wysiwyg = "true";
defparam \mem[50][67] .power_up = "low";

cycloneive_lcell_comb \mem[49][67]~98 (
	.dataa(\mem[50][67]~q ),
	.datab(\mem_used[50]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[49][67]~98_combout ),
	.cout());
defparam \mem[49][67]~98 .lut_mask = 16'hB8FF;
defparam \mem[49][67]~98 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[49][67]~99 (
	.dataa(\mem[49][67]~q ),
	.datab(\mem[49][67]~98_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[49]~q ),
	.cin(gnd),
	.combout(\mem[49][67]~99_combout ),
	.cout());
defparam \mem[49][67]~99 .lut_mask = 16'hEFFE;
defparam \mem[49][67]~99 .sum_lutc_input = "datac";

dffeas \mem[49][67] (
	.clk(clk),
	.d(\mem[49][67]~99_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[49][67]~q ),
	.prn(vcc));
defparam \mem[49][67] .is_wysiwyg = "true";
defparam \mem[49][67] .power_up = "low";

cycloneive_lcell_comb \mem[48][67]~96 (
	.dataa(\mem[49][67]~q ),
	.datab(\mem_used[49]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[48][67]~96_combout ),
	.cout());
defparam \mem[48][67]~96 .lut_mask = 16'hB8FF;
defparam \mem[48][67]~96 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[48][67]~97 (
	.dataa(\mem[48][67]~q ),
	.datab(\mem[48][67]~96_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[48]~q ),
	.cin(gnd),
	.combout(\mem[48][67]~97_combout ),
	.cout());
defparam \mem[48][67]~97 .lut_mask = 16'hEFFE;
defparam \mem[48][67]~97 .sum_lutc_input = "datac";

dffeas \mem[48][67] (
	.clk(clk),
	.d(\mem[48][67]~97_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[48][67]~q ),
	.prn(vcc));
defparam \mem[48][67] .is_wysiwyg = "true";
defparam \mem[48][67] .power_up = "low";

cycloneive_lcell_comb \mem[47][67]~94 (
	.dataa(\mem[48][67]~q ),
	.datab(\mem_used[48]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[47][67]~94_combout ),
	.cout());
defparam \mem[47][67]~94 .lut_mask = 16'hB8FF;
defparam \mem[47][67]~94 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[47][67]~95 (
	.dataa(\mem[47][67]~q ),
	.datab(\mem[47][67]~94_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[47]~q ),
	.cin(gnd),
	.combout(\mem[47][67]~95_combout ),
	.cout());
defparam \mem[47][67]~95 .lut_mask = 16'hEFFE;
defparam \mem[47][67]~95 .sum_lutc_input = "datac";

dffeas \mem[47][67] (
	.clk(clk),
	.d(\mem[47][67]~95_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[47][67]~q ),
	.prn(vcc));
defparam \mem[47][67] .is_wysiwyg = "true";
defparam \mem[47][67] .power_up = "low";

cycloneive_lcell_comb \mem[46][67]~92 (
	.dataa(\mem[47][67]~q ),
	.datab(\mem_used[47]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[46][67]~92_combout ),
	.cout());
defparam \mem[46][67]~92 .lut_mask = 16'hB8FF;
defparam \mem[46][67]~92 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[46][67]~93 (
	.dataa(\mem[46][67]~q ),
	.datab(\mem[46][67]~92_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[46]~q ),
	.cin(gnd),
	.combout(\mem[46][67]~93_combout ),
	.cout());
defparam \mem[46][67]~93 .lut_mask = 16'hEFFE;
defparam \mem[46][67]~93 .sum_lutc_input = "datac";

dffeas \mem[46][67] (
	.clk(clk),
	.d(\mem[46][67]~93_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[46][67]~q ),
	.prn(vcc));
defparam \mem[46][67] .is_wysiwyg = "true";
defparam \mem[46][67] .power_up = "low";

cycloneive_lcell_comb \mem[45][67]~90 (
	.dataa(\mem[46][67]~q ),
	.datab(\mem_used[46]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[45][67]~90_combout ),
	.cout());
defparam \mem[45][67]~90 .lut_mask = 16'hB8FF;
defparam \mem[45][67]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[45][67]~91 (
	.dataa(\mem[45][67]~q ),
	.datab(\mem[45][67]~90_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[45]~q ),
	.cin(gnd),
	.combout(\mem[45][67]~91_combout ),
	.cout());
defparam \mem[45][67]~91 .lut_mask = 16'hEFFE;
defparam \mem[45][67]~91 .sum_lutc_input = "datac";

dffeas \mem[45][67] (
	.clk(clk),
	.d(\mem[45][67]~91_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[45][67]~q ),
	.prn(vcc));
defparam \mem[45][67] .is_wysiwyg = "true";
defparam \mem[45][67] .power_up = "low";

cycloneive_lcell_comb \mem[44][67]~88 (
	.dataa(\mem[45][67]~q ),
	.datab(\mem_used[45]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[44][67]~88_combout ),
	.cout());
defparam \mem[44][67]~88 .lut_mask = 16'hB8FF;
defparam \mem[44][67]~88 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[44][67]~89 (
	.dataa(\mem[44][67]~q ),
	.datab(\mem[44][67]~88_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[44]~q ),
	.cin(gnd),
	.combout(\mem[44][67]~89_combout ),
	.cout());
defparam \mem[44][67]~89 .lut_mask = 16'hEFFE;
defparam \mem[44][67]~89 .sum_lutc_input = "datac";

dffeas \mem[44][67] (
	.clk(clk),
	.d(\mem[44][67]~89_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[44][67]~q ),
	.prn(vcc));
defparam \mem[44][67] .is_wysiwyg = "true";
defparam \mem[44][67] .power_up = "low";

cycloneive_lcell_comb \mem[43][67]~86 (
	.dataa(\mem[44][67]~q ),
	.datab(\mem_used[44]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[43][67]~86_combout ),
	.cout());
defparam \mem[43][67]~86 .lut_mask = 16'hB8FF;
defparam \mem[43][67]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[43][67]~87 (
	.dataa(\mem[43][67]~q ),
	.datab(\mem[43][67]~86_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[43]~q ),
	.cin(gnd),
	.combout(\mem[43][67]~87_combout ),
	.cout());
defparam \mem[43][67]~87 .lut_mask = 16'hEFFE;
defparam \mem[43][67]~87 .sum_lutc_input = "datac";

dffeas \mem[43][67] (
	.clk(clk),
	.d(\mem[43][67]~87_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[43][67]~q ),
	.prn(vcc));
defparam \mem[43][67] .is_wysiwyg = "true";
defparam \mem[43][67] .power_up = "low";

cycloneive_lcell_comb \mem[42][67]~84 (
	.dataa(\mem[43][67]~q ),
	.datab(\mem_used[43]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[42][67]~84_combout ),
	.cout());
defparam \mem[42][67]~84 .lut_mask = 16'hB8FF;
defparam \mem[42][67]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[42][67]~85 (
	.dataa(\mem[42][67]~q ),
	.datab(\mem[42][67]~84_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[42]~q ),
	.cin(gnd),
	.combout(\mem[42][67]~85_combout ),
	.cout());
defparam \mem[42][67]~85 .lut_mask = 16'hEFFE;
defparam \mem[42][67]~85 .sum_lutc_input = "datac";

dffeas \mem[42][67] (
	.clk(clk),
	.d(\mem[42][67]~85_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[42][67]~q ),
	.prn(vcc));
defparam \mem[42][67] .is_wysiwyg = "true";
defparam \mem[42][67] .power_up = "low";

cycloneive_lcell_comb \mem[41][67]~82 (
	.dataa(\mem[42][67]~q ),
	.datab(\mem_used[42]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[41][67]~82_combout ),
	.cout());
defparam \mem[41][67]~82 .lut_mask = 16'hB8FF;
defparam \mem[41][67]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[41][67]~83 (
	.dataa(\mem[41][67]~q ),
	.datab(\mem[41][67]~82_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[41]~q ),
	.cin(gnd),
	.combout(\mem[41][67]~83_combout ),
	.cout());
defparam \mem[41][67]~83 .lut_mask = 16'hEFFE;
defparam \mem[41][67]~83 .sum_lutc_input = "datac";

dffeas \mem[41][67] (
	.clk(clk),
	.d(\mem[41][67]~83_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[41][67]~q ),
	.prn(vcc));
defparam \mem[41][67] .is_wysiwyg = "true";
defparam \mem[41][67] .power_up = "low";

cycloneive_lcell_comb \mem[40][67]~80 (
	.dataa(\mem[41][67]~q ),
	.datab(\mem_used[41]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[40][67]~80_combout ),
	.cout());
defparam \mem[40][67]~80 .lut_mask = 16'hB8FF;
defparam \mem[40][67]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[40][67]~81 (
	.dataa(\mem[40][67]~q ),
	.datab(\mem[40][67]~80_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[40]~q ),
	.cin(gnd),
	.combout(\mem[40][67]~81_combout ),
	.cout());
defparam \mem[40][67]~81 .lut_mask = 16'hEFFE;
defparam \mem[40][67]~81 .sum_lutc_input = "datac";

dffeas \mem[40][67] (
	.clk(clk),
	.d(\mem[40][67]~81_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[40][67]~q ),
	.prn(vcc));
defparam \mem[40][67] .is_wysiwyg = "true";
defparam \mem[40][67] .power_up = "low";

cycloneive_lcell_comb \mem[39][67]~78 (
	.dataa(\mem[40][67]~q ),
	.datab(\mem_used[40]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[39][67]~78_combout ),
	.cout());
defparam \mem[39][67]~78 .lut_mask = 16'hB8FF;
defparam \mem[39][67]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[39][67]~79 (
	.dataa(\mem[39][67]~q ),
	.datab(\mem[39][67]~78_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[39]~q ),
	.cin(gnd),
	.combout(\mem[39][67]~79_combout ),
	.cout());
defparam \mem[39][67]~79 .lut_mask = 16'hEFFE;
defparam \mem[39][67]~79 .sum_lutc_input = "datac";

dffeas \mem[39][67] (
	.clk(clk),
	.d(\mem[39][67]~79_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[39][67]~q ),
	.prn(vcc));
defparam \mem[39][67] .is_wysiwyg = "true";
defparam \mem[39][67] .power_up = "low";

cycloneive_lcell_comb \mem[38][67]~76 (
	.dataa(\mem[39][67]~q ),
	.datab(\mem_used[39]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[38][67]~76_combout ),
	.cout());
defparam \mem[38][67]~76 .lut_mask = 16'hB8FF;
defparam \mem[38][67]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[38][67]~77 (
	.dataa(\mem[38][67]~q ),
	.datab(\mem[38][67]~76_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[38]~q ),
	.cin(gnd),
	.combout(\mem[38][67]~77_combout ),
	.cout());
defparam \mem[38][67]~77 .lut_mask = 16'hEFFE;
defparam \mem[38][67]~77 .sum_lutc_input = "datac";

dffeas \mem[38][67] (
	.clk(clk),
	.d(\mem[38][67]~77_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[38][67]~q ),
	.prn(vcc));
defparam \mem[38][67] .is_wysiwyg = "true";
defparam \mem[38][67] .power_up = "low";

cycloneive_lcell_comb \mem[37][67]~74 (
	.dataa(\mem[38][67]~q ),
	.datab(\mem_used[38]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[37][67]~74_combout ),
	.cout());
defparam \mem[37][67]~74 .lut_mask = 16'hB8FF;
defparam \mem[37][67]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[37][67]~75 (
	.dataa(\mem[37][67]~q ),
	.datab(\mem[37][67]~74_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[37]~q ),
	.cin(gnd),
	.combout(\mem[37][67]~75_combout ),
	.cout());
defparam \mem[37][67]~75 .lut_mask = 16'hEFFE;
defparam \mem[37][67]~75 .sum_lutc_input = "datac";

dffeas \mem[37][67] (
	.clk(clk),
	.d(\mem[37][67]~75_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[37][67]~q ),
	.prn(vcc));
defparam \mem[37][67] .is_wysiwyg = "true";
defparam \mem[37][67] .power_up = "low";

cycloneive_lcell_comb \mem[36][67]~72 (
	.dataa(\mem[37][67]~q ),
	.datab(\mem_used[37]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[36][67]~72_combout ),
	.cout());
defparam \mem[36][67]~72 .lut_mask = 16'hB8FF;
defparam \mem[36][67]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[36][67]~73 (
	.dataa(\mem[36][67]~q ),
	.datab(\mem[36][67]~72_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[36]~q ),
	.cin(gnd),
	.combout(\mem[36][67]~73_combout ),
	.cout());
defparam \mem[36][67]~73 .lut_mask = 16'hEFFE;
defparam \mem[36][67]~73 .sum_lutc_input = "datac";

dffeas \mem[36][67] (
	.clk(clk),
	.d(\mem[36][67]~73_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[36][67]~q ),
	.prn(vcc));
defparam \mem[36][67] .is_wysiwyg = "true";
defparam \mem[36][67] .power_up = "low";

cycloneive_lcell_comb \mem[35][67]~70 (
	.dataa(\mem[36][67]~q ),
	.datab(\mem_used[36]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[35][67]~70_combout ),
	.cout());
defparam \mem[35][67]~70 .lut_mask = 16'hB8FF;
defparam \mem[35][67]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[35][67]~71 (
	.dataa(\mem[35][67]~q ),
	.datab(\mem[35][67]~70_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[35]~q ),
	.cin(gnd),
	.combout(\mem[35][67]~71_combout ),
	.cout());
defparam \mem[35][67]~71 .lut_mask = 16'hEFFE;
defparam \mem[35][67]~71 .sum_lutc_input = "datac";

dffeas \mem[35][67] (
	.clk(clk),
	.d(\mem[35][67]~71_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[35][67]~q ),
	.prn(vcc));
defparam \mem[35][67] .is_wysiwyg = "true";
defparam \mem[35][67] .power_up = "low";

cycloneive_lcell_comb \mem[34][67]~68 (
	.dataa(\mem[35][67]~q ),
	.datab(\mem_used[35]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[34][67]~68_combout ),
	.cout());
defparam \mem[34][67]~68 .lut_mask = 16'hB8FF;
defparam \mem[34][67]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[34][67]~69 (
	.dataa(\mem[34][67]~q ),
	.datab(\mem[34][67]~68_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[34]~q ),
	.cin(gnd),
	.combout(\mem[34][67]~69_combout ),
	.cout());
defparam \mem[34][67]~69 .lut_mask = 16'hEFFE;
defparam \mem[34][67]~69 .sum_lutc_input = "datac";

dffeas \mem[34][67] (
	.clk(clk),
	.d(\mem[34][67]~69_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[34][67]~q ),
	.prn(vcc));
defparam \mem[34][67] .is_wysiwyg = "true";
defparam \mem[34][67] .power_up = "low";

cycloneive_lcell_comb \mem[33][67]~66 (
	.dataa(\mem[34][67]~q ),
	.datab(\mem_used[34]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[33][67]~66_combout ),
	.cout());
defparam \mem[33][67]~66 .lut_mask = 16'hB8FF;
defparam \mem[33][67]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[33][67]~67 (
	.dataa(\mem[33][67]~q ),
	.datab(\mem[33][67]~66_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[33]~q ),
	.cin(gnd),
	.combout(\mem[33][67]~67_combout ),
	.cout());
defparam \mem[33][67]~67 .lut_mask = 16'hEFFE;
defparam \mem[33][67]~67 .sum_lutc_input = "datac";

dffeas \mem[33][67] (
	.clk(clk),
	.d(\mem[33][67]~67_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[33][67]~q ),
	.prn(vcc));
defparam \mem[33][67] .is_wysiwyg = "true";
defparam \mem[33][67] .power_up = "low";

cycloneive_lcell_comb \mem[32][67]~64 (
	.dataa(\mem[33][67]~q ),
	.datab(\mem_used[33]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[32][67]~64_combout ),
	.cout());
defparam \mem[32][67]~64 .lut_mask = 16'hB8FF;
defparam \mem[32][67]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[32][67]~65 (
	.dataa(\mem[32][67]~q ),
	.datab(\mem[32][67]~64_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[32]~q ),
	.cin(gnd),
	.combout(\mem[32][67]~65_combout ),
	.cout());
defparam \mem[32][67]~65 .lut_mask = 16'hEFFE;
defparam \mem[32][67]~65 .sum_lutc_input = "datac";

dffeas \mem[32][67] (
	.clk(clk),
	.d(\mem[32][67]~65_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[32][67]~q ),
	.prn(vcc));
defparam \mem[32][67] .is_wysiwyg = "true";
defparam \mem[32][67] .power_up = "low";

cycloneive_lcell_comb \mem[31][67]~62 (
	.dataa(\mem[32][67]~q ),
	.datab(\mem_used[32]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[31][67]~62_combout ),
	.cout());
defparam \mem[31][67]~62 .lut_mask = 16'hB8FF;
defparam \mem[31][67]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[31][67]~63 (
	.dataa(\mem[31][67]~q ),
	.datab(\mem[31][67]~62_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[31]~q ),
	.cin(gnd),
	.combout(\mem[31][67]~63_combout ),
	.cout());
defparam \mem[31][67]~63 .lut_mask = 16'hEFFE;
defparam \mem[31][67]~63 .sum_lutc_input = "datac";

dffeas \mem[31][67] (
	.clk(clk),
	.d(\mem[31][67]~63_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[31][67]~q ),
	.prn(vcc));
defparam \mem[31][67] .is_wysiwyg = "true";
defparam \mem[31][67] .power_up = "low";

cycloneive_lcell_comb \mem[30][67]~60 (
	.dataa(\mem[31][67]~q ),
	.datab(\mem_used[31]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[30][67]~60_combout ),
	.cout());
defparam \mem[30][67]~60 .lut_mask = 16'hB8FF;
defparam \mem[30][67]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[30][67]~61 (
	.dataa(\mem[30][67]~q ),
	.datab(\mem[30][67]~60_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[30]~q ),
	.cin(gnd),
	.combout(\mem[30][67]~61_combout ),
	.cout());
defparam \mem[30][67]~61 .lut_mask = 16'hEFFE;
defparam \mem[30][67]~61 .sum_lutc_input = "datac";

dffeas \mem[30][67] (
	.clk(clk),
	.d(\mem[30][67]~61_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[30][67]~q ),
	.prn(vcc));
defparam \mem[30][67] .is_wysiwyg = "true";
defparam \mem[30][67] .power_up = "low";

cycloneive_lcell_comb \mem[29][67]~58 (
	.dataa(\mem[30][67]~q ),
	.datab(\mem_used[30]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[29][67]~58_combout ),
	.cout());
defparam \mem[29][67]~58 .lut_mask = 16'hB8FF;
defparam \mem[29][67]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[29][67]~59 (
	.dataa(\mem[29][67]~q ),
	.datab(\mem[29][67]~58_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[29]~q ),
	.cin(gnd),
	.combout(\mem[29][67]~59_combout ),
	.cout());
defparam \mem[29][67]~59 .lut_mask = 16'hEFFE;
defparam \mem[29][67]~59 .sum_lutc_input = "datac";

dffeas \mem[29][67] (
	.clk(clk),
	.d(\mem[29][67]~59_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[29][67]~q ),
	.prn(vcc));
defparam \mem[29][67] .is_wysiwyg = "true";
defparam \mem[29][67] .power_up = "low";

cycloneive_lcell_comb \mem[28][67]~56 (
	.dataa(\mem[29][67]~q ),
	.datab(\mem_used[29]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[28][67]~56_combout ),
	.cout());
defparam \mem[28][67]~56 .lut_mask = 16'hB8FF;
defparam \mem[28][67]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[28][67]~57 (
	.dataa(\mem[28][67]~q ),
	.datab(\mem[28][67]~56_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[28]~q ),
	.cin(gnd),
	.combout(\mem[28][67]~57_combout ),
	.cout());
defparam \mem[28][67]~57 .lut_mask = 16'hEFFE;
defparam \mem[28][67]~57 .sum_lutc_input = "datac";

dffeas \mem[28][67] (
	.clk(clk),
	.d(\mem[28][67]~57_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[28][67]~q ),
	.prn(vcc));
defparam \mem[28][67] .is_wysiwyg = "true";
defparam \mem[28][67] .power_up = "low";

cycloneive_lcell_comb \mem[27][67]~54 (
	.dataa(\mem[28][67]~q ),
	.datab(\mem_used[28]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[27][67]~54_combout ),
	.cout());
defparam \mem[27][67]~54 .lut_mask = 16'hB8FF;
defparam \mem[27][67]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[27][67]~55 (
	.dataa(\mem[27][67]~q ),
	.datab(\mem[27][67]~54_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[27]~q ),
	.cin(gnd),
	.combout(\mem[27][67]~55_combout ),
	.cout());
defparam \mem[27][67]~55 .lut_mask = 16'hEFFE;
defparam \mem[27][67]~55 .sum_lutc_input = "datac";

dffeas \mem[27][67] (
	.clk(clk),
	.d(\mem[27][67]~55_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[27][67]~q ),
	.prn(vcc));
defparam \mem[27][67] .is_wysiwyg = "true";
defparam \mem[27][67] .power_up = "low";

cycloneive_lcell_comb \mem[26][67]~52 (
	.dataa(\mem[27][67]~q ),
	.datab(\mem_used[27]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[26][67]~52_combout ),
	.cout());
defparam \mem[26][67]~52 .lut_mask = 16'hB8FF;
defparam \mem[26][67]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[26][67]~53 (
	.dataa(\mem[26][67]~q ),
	.datab(\mem[26][67]~52_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[26]~q ),
	.cin(gnd),
	.combout(\mem[26][67]~53_combout ),
	.cout());
defparam \mem[26][67]~53 .lut_mask = 16'hEFFE;
defparam \mem[26][67]~53 .sum_lutc_input = "datac";

dffeas \mem[26][67] (
	.clk(clk),
	.d(\mem[26][67]~53_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[26][67]~q ),
	.prn(vcc));
defparam \mem[26][67] .is_wysiwyg = "true";
defparam \mem[26][67] .power_up = "low";

cycloneive_lcell_comb \mem[25][67]~50 (
	.dataa(\mem[26][67]~q ),
	.datab(\mem_used[26]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[25][67]~50_combout ),
	.cout());
defparam \mem[25][67]~50 .lut_mask = 16'hB8FF;
defparam \mem[25][67]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[25][67]~51 (
	.dataa(\mem[25][67]~q ),
	.datab(\mem[25][67]~50_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[25]~q ),
	.cin(gnd),
	.combout(\mem[25][67]~51_combout ),
	.cout());
defparam \mem[25][67]~51 .lut_mask = 16'hEFFE;
defparam \mem[25][67]~51 .sum_lutc_input = "datac";

dffeas \mem[25][67] (
	.clk(clk),
	.d(\mem[25][67]~51_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[25][67]~q ),
	.prn(vcc));
defparam \mem[25][67] .is_wysiwyg = "true";
defparam \mem[25][67] .power_up = "low";

cycloneive_lcell_comb \mem[24][67]~48 (
	.dataa(\mem[25][67]~q ),
	.datab(\mem_used[25]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[24][67]~48_combout ),
	.cout());
defparam \mem[24][67]~48 .lut_mask = 16'hB8FF;
defparam \mem[24][67]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[24][67]~49 (
	.dataa(\mem[24][67]~q ),
	.datab(\mem[24][67]~48_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[24]~q ),
	.cin(gnd),
	.combout(\mem[24][67]~49_combout ),
	.cout());
defparam \mem[24][67]~49 .lut_mask = 16'hEFFE;
defparam \mem[24][67]~49 .sum_lutc_input = "datac";

dffeas \mem[24][67] (
	.clk(clk),
	.d(\mem[24][67]~49_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[24][67]~q ),
	.prn(vcc));
defparam \mem[24][67] .is_wysiwyg = "true";
defparam \mem[24][67] .power_up = "low";

cycloneive_lcell_comb \mem[23][67]~46 (
	.dataa(\mem[24][67]~q ),
	.datab(\mem_used[24]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[23][67]~46_combout ),
	.cout());
defparam \mem[23][67]~46 .lut_mask = 16'hB8FF;
defparam \mem[23][67]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[23][67]~47 (
	.dataa(\mem[23][67]~q ),
	.datab(\mem[23][67]~46_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[23]~q ),
	.cin(gnd),
	.combout(\mem[23][67]~47_combout ),
	.cout());
defparam \mem[23][67]~47 .lut_mask = 16'hEFFE;
defparam \mem[23][67]~47 .sum_lutc_input = "datac";

dffeas \mem[23][67] (
	.clk(clk),
	.d(\mem[23][67]~47_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[23][67]~q ),
	.prn(vcc));
defparam \mem[23][67] .is_wysiwyg = "true";
defparam \mem[23][67] .power_up = "low";

cycloneive_lcell_comb \mem[22][67]~44 (
	.dataa(\mem[23][67]~q ),
	.datab(\mem_used[23]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[22][67]~44_combout ),
	.cout());
defparam \mem[22][67]~44 .lut_mask = 16'hB8FF;
defparam \mem[22][67]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[22][67]~45 (
	.dataa(\mem[22][67]~q ),
	.datab(\mem[22][67]~44_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[22]~q ),
	.cin(gnd),
	.combout(\mem[22][67]~45_combout ),
	.cout());
defparam \mem[22][67]~45 .lut_mask = 16'hEFFE;
defparam \mem[22][67]~45 .sum_lutc_input = "datac";

dffeas \mem[22][67] (
	.clk(clk),
	.d(\mem[22][67]~45_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[22][67]~q ),
	.prn(vcc));
defparam \mem[22][67] .is_wysiwyg = "true";
defparam \mem[22][67] .power_up = "low";

cycloneive_lcell_comb \mem[21][67]~42 (
	.dataa(\mem[22][67]~q ),
	.datab(\mem_used[22]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[21][67]~42_combout ),
	.cout());
defparam \mem[21][67]~42 .lut_mask = 16'hB8FF;
defparam \mem[21][67]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[21][67]~43 (
	.dataa(\mem[21][67]~q ),
	.datab(\mem[21][67]~42_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[21]~q ),
	.cin(gnd),
	.combout(\mem[21][67]~43_combout ),
	.cout());
defparam \mem[21][67]~43 .lut_mask = 16'hEFFE;
defparam \mem[21][67]~43 .sum_lutc_input = "datac";

dffeas \mem[21][67] (
	.clk(clk),
	.d(\mem[21][67]~43_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[21][67]~q ),
	.prn(vcc));
defparam \mem[21][67] .is_wysiwyg = "true";
defparam \mem[21][67] .power_up = "low";

cycloneive_lcell_comb \mem[20][67]~40 (
	.dataa(\mem[21][67]~q ),
	.datab(\mem_used[21]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[20][67]~40_combout ),
	.cout());
defparam \mem[20][67]~40 .lut_mask = 16'hB8FF;
defparam \mem[20][67]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[20][67]~41 (
	.dataa(\mem[20][67]~q ),
	.datab(\mem[20][67]~40_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[20]~q ),
	.cin(gnd),
	.combout(\mem[20][67]~41_combout ),
	.cout());
defparam \mem[20][67]~41 .lut_mask = 16'hEFFE;
defparam \mem[20][67]~41 .sum_lutc_input = "datac";

dffeas \mem[20][67] (
	.clk(clk),
	.d(\mem[20][67]~41_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[20][67]~q ),
	.prn(vcc));
defparam \mem[20][67] .is_wysiwyg = "true";
defparam \mem[20][67] .power_up = "low";

cycloneive_lcell_comb \mem[19][67]~38 (
	.dataa(\mem[20][67]~q ),
	.datab(\mem_used[20]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[19][67]~38_combout ),
	.cout());
defparam \mem[19][67]~38 .lut_mask = 16'hB8FF;
defparam \mem[19][67]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[19][67]~39 (
	.dataa(\mem[19][67]~q ),
	.datab(\mem[19][67]~38_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[19]~q ),
	.cin(gnd),
	.combout(\mem[19][67]~39_combout ),
	.cout());
defparam \mem[19][67]~39 .lut_mask = 16'hEFFE;
defparam \mem[19][67]~39 .sum_lutc_input = "datac";

dffeas \mem[19][67] (
	.clk(clk),
	.d(\mem[19][67]~39_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[19][67]~q ),
	.prn(vcc));
defparam \mem[19][67] .is_wysiwyg = "true";
defparam \mem[19][67] .power_up = "low";

cycloneive_lcell_comb \mem[18][67]~36 (
	.dataa(\mem[19][67]~q ),
	.datab(\mem_used[19]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[18][67]~36_combout ),
	.cout());
defparam \mem[18][67]~36 .lut_mask = 16'hB8FF;
defparam \mem[18][67]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[18][67]~37 (
	.dataa(\mem[18][67]~q ),
	.datab(\mem[18][67]~36_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[18]~q ),
	.cin(gnd),
	.combout(\mem[18][67]~37_combout ),
	.cout());
defparam \mem[18][67]~37 .lut_mask = 16'hEFFE;
defparam \mem[18][67]~37 .sum_lutc_input = "datac";

dffeas \mem[18][67] (
	.clk(clk),
	.d(\mem[18][67]~37_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[18][67]~q ),
	.prn(vcc));
defparam \mem[18][67] .is_wysiwyg = "true";
defparam \mem[18][67] .power_up = "low";

cycloneive_lcell_comb \mem[17][67]~34 (
	.dataa(\mem[18][67]~q ),
	.datab(\mem_used[18]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[17][67]~34_combout ),
	.cout());
defparam \mem[17][67]~34 .lut_mask = 16'hB8FF;
defparam \mem[17][67]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[17][67]~35 (
	.dataa(\mem[17][67]~q ),
	.datab(\mem[17][67]~34_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[17]~q ),
	.cin(gnd),
	.combout(\mem[17][67]~35_combout ),
	.cout());
defparam \mem[17][67]~35 .lut_mask = 16'hEFFE;
defparam \mem[17][67]~35 .sum_lutc_input = "datac";

dffeas \mem[17][67] (
	.clk(clk),
	.d(\mem[17][67]~35_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[17][67]~q ),
	.prn(vcc));
defparam \mem[17][67] .is_wysiwyg = "true";
defparam \mem[17][67] .power_up = "low";

cycloneive_lcell_comb \mem[16][67]~32 (
	.dataa(\mem[17][67]~q ),
	.datab(\mem_used[17]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[16][67]~32_combout ),
	.cout());
defparam \mem[16][67]~32 .lut_mask = 16'hB8FF;
defparam \mem[16][67]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[16][67]~33 (
	.dataa(\mem[16][67]~q ),
	.datab(\mem[16][67]~32_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[16]~q ),
	.cin(gnd),
	.combout(\mem[16][67]~33_combout ),
	.cout());
defparam \mem[16][67]~33 .lut_mask = 16'hEFFE;
defparam \mem[16][67]~33 .sum_lutc_input = "datac";

dffeas \mem[16][67] (
	.clk(clk),
	.d(\mem[16][67]~33_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[16][67]~q ),
	.prn(vcc));
defparam \mem[16][67] .is_wysiwyg = "true";
defparam \mem[16][67] .power_up = "low";

cycloneive_lcell_comb \mem[15][67]~30 (
	.dataa(\mem[16][67]~q ),
	.datab(\mem_used[16]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[15][67]~30_combout ),
	.cout());
defparam \mem[15][67]~30 .lut_mask = 16'hB8FF;
defparam \mem[15][67]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[15][67]~31 (
	.dataa(\mem[15][67]~q ),
	.datab(\mem[15][67]~30_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[15]~q ),
	.cin(gnd),
	.combout(\mem[15][67]~31_combout ),
	.cout());
defparam \mem[15][67]~31 .lut_mask = 16'hEFFE;
defparam \mem[15][67]~31 .sum_lutc_input = "datac";

dffeas \mem[15][67] (
	.clk(clk),
	.d(\mem[15][67]~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[15][67]~q ),
	.prn(vcc));
defparam \mem[15][67] .is_wysiwyg = "true";
defparam \mem[15][67] .power_up = "low";

cycloneive_lcell_comb \mem[14][67]~28 (
	.dataa(\mem[15][67]~q ),
	.datab(\mem_used[15]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[14][67]~28_combout ),
	.cout());
defparam \mem[14][67]~28 .lut_mask = 16'hB8FF;
defparam \mem[14][67]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[14][67]~29 (
	.dataa(\mem[14][67]~q ),
	.datab(\mem[14][67]~28_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[14]~q ),
	.cin(gnd),
	.combout(\mem[14][67]~29_combout ),
	.cout());
defparam \mem[14][67]~29 .lut_mask = 16'hEFFE;
defparam \mem[14][67]~29 .sum_lutc_input = "datac";

dffeas \mem[14][67] (
	.clk(clk),
	.d(\mem[14][67]~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[14][67]~q ),
	.prn(vcc));
defparam \mem[14][67] .is_wysiwyg = "true";
defparam \mem[14][67] .power_up = "low";

cycloneive_lcell_comb \mem[13][67]~26 (
	.dataa(\mem[14][67]~q ),
	.datab(\mem_used[14]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[13][67]~26_combout ),
	.cout());
defparam \mem[13][67]~26 .lut_mask = 16'hB8FF;
defparam \mem[13][67]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[13][67]~27 (
	.dataa(\mem[13][67]~q ),
	.datab(\mem[13][67]~26_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[13]~q ),
	.cin(gnd),
	.combout(\mem[13][67]~27_combout ),
	.cout());
defparam \mem[13][67]~27 .lut_mask = 16'hEFFE;
defparam \mem[13][67]~27 .sum_lutc_input = "datac";

dffeas \mem[13][67] (
	.clk(clk),
	.d(\mem[13][67]~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[13][67]~q ),
	.prn(vcc));
defparam \mem[13][67] .is_wysiwyg = "true";
defparam \mem[13][67] .power_up = "low";

cycloneive_lcell_comb \mem[12][67]~24 (
	.dataa(\mem[13][67]~q ),
	.datab(\mem_used[13]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[12][67]~24_combout ),
	.cout());
defparam \mem[12][67]~24 .lut_mask = 16'hB8FF;
defparam \mem[12][67]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[12][67]~25 (
	.dataa(\mem[12][67]~q ),
	.datab(\mem[12][67]~24_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[12]~q ),
	.cin(gnd),
	.combout(\mem[12][67]~25_combout ),
	.cout());
defparam \mem[12][67]~25 .lut_mask = 16'hEFFE;
defparam \mem[12][67]~25 .sum_lutc_input = "datac";

dffeas \mem[12][67] (
	.clk(clk),
	.d(\mem[12][67]~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[12][67]~q ),
	.prn(vcc));
defparam \mem[12][67] .is_wysiwyg = "true";
defparam \mem[12][67] .power_up = "low";

cycloneive_lcell_comb \mem[11][67]~22 (
	.dataa(\mem[12][67]~q ),
	.datab(\mem_used[12]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[11][67]~22_combout ),
	.cout());
defparam \mem[11][67]~22 .lut_mask = 16'hB8FF;
defparam \mem[11][67]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[11][67]~23 (
	.dataa(\mem[11][67]~q ),
	.datab(\mem[11][67]~22_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[11]~q ),
	.cin(gnd),
	.combout(\mem[11][67]~23_combout ),
	.cout());
defparam \mem[11][67]~23 .lut_mask = 16'hEFFE;
defparam \mem[11][67]~23 .sum_lutc_input = "datac";

dffeas \mem[11][67] (
	.clk(clk),
	.d(\mem[11][67]~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[11][67]~q ),
	.prn(vcc));
defparam \mem[11][67] .is_wysiwyg = "true";
defparam \mem[11][67] .power_up = "low";

cycloneive_lcell_comb \mem[10][67]~20 (
	.dataa(\mem[11][67]~q ),
	.datab(\mem_used[11]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[10][67]~20_combout ),
	.cout());
defparam \mem[10][67]~20 .lut_mask = 16'hB8FF;
defparam \mem[10][67]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[10][67]~21 (
	.dataa(\mem[10][67]~q ),
	.datab(\mem[10][67]~20_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[10]~q ),
	.cin(gnd),
	.combout(\mem[10][67]~21_combout ),
	.cout());
defparam \mem[10][67]~21 .lut_mask = 16'hEFFE;
defparam \mem[10][67]~21 .sum_lutc_input = "datac";

dffeas \mem[10][67] (
	.clk(clk),
	.d(\mem[10][67]~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[10][67]~q ),
	.prn(vcc));
defparam \mem[10][67] .is_wysiwyg = "true";
defparam \mem[10][67] .power_up = "low";

cycloneive_lcell_comb \mem[9][67]~18 (
	.dataa(\mem[10][67]~q ),
	.datab(\mem_used[10]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[9][67]~18_combout ),
	.cout());
defparam \mem[9][67]~18 .lut_mask = 16'hB8FF;
defparam \mem[9][67]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[9][67]~19 (
	.dataa(\mem[9][67]~q ),
	.datab(\mem[9][67]~18_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[9]~q ),
	.cin(gnd),
	.combout(\mem[9][67]~19_combout ),
	.cout());
defparam \mem[9][67]~19 .lut_mask = 16'hEFFE;
defparam \mem[9][67]~19 .sum_lutc_input = "datac";

dffeas \mem[9][67] (
	.clk(clk),
	.d(\mem[9][67]~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][67]~q ),
	.prn(vcc));
defparam \mem[9][67] .is_wysiwyg = "true";
defparam \mem[9][67] .power_up = "low";

cycloneive_lcell_comb \mem[8][67]~16 (
	.dataa(\mem[9][67]~q ),
	.datab(\mem_used[9]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[8][67]~16_combout ),
	.cout());
defparam \mem[8][67]~16 .lut_mask = 16'hB8FF;
defparam \mem[8][67]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[8][67]~17 (
	.dataa(\mem[8][67]~q ),
	.datab(\mem[8][67]~16_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem[8][67]~17_combout ),
	.cout());
defparam \mem[8][67]~17 .lut_mask = 16'hEFFE;
defparam \mem[8][67]~17 .sum_lutc_input = "datac";

dffeas \mem[8][67] (
	.clk(clk),
	.d(\mem[8][67]~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[8][67]~q ),
	.prn(vcc));
defparam \mem[8][67] .is_wysiwyg = "true";
defparam \mem[8][67] .power_up = "low";

cycloneive_lcell_comb \mem[7][67]~14 (
	.dataa(\mem[8][67]~q ),
	.datab(\mem_used[8]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[7][67]~14_combout ),
	.cout());
defparam \mem[7][67]~14 .lut_mask = 16'hB8FF;
defparam \mem[7][67]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[7][67]~15 (
	.dataa(\mem[7][67]~q ),
	.datab(\mem[7][67]~14_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem[7][67]~15_combout ),
	.cout());
defparam \mem[7][67]~15 .lut_mask = 16'hEFFE;
defparam \mem[7][67]~15 .sum_lutc_input = "datac";

dffeas \mem[7][67] (
	.clk(clk),
	.d(\mem[7][67]~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][67]~q ),
	.prn(vcc));
defparam \mem[7][67] .is_wysiwyg = "true";
defparam \mem[7][67] .power_up = "low";

cycloneive_lcell_comb \mem[6][67]~12 (
	.dataa(\mem[7][67]~q ),
	.datab(\mem_used[7]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[6][67]~12_combout ),
	.cout());
defparam \mem[6][67]~12 .lut_mask = 16'hB8FF;
defparam \mem[6][67]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[6][67]~13 (
	.dataa(\mem[6][67]~q ),
	.datab(\mem[6][67]~12_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem[6][67]~13_combout ),
	.cout());
defparam \mem[6][67]~13 .lut_mask = 16'hEFFE;
defparam \mem[6][67]~13 .sum_lutc_input = "datac";

dffeas \mem[6][67] (
	.clk(clk),
	.d(\mem[6][67]~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[6][67]~q ),
	.prn(vcc));
defparam \mem[6][67] .is_wysiwyg = "true";
defparam \mem[6][67] .power_up = "low";

cycloneive_lcell_comb \mem[5][67]~10 (
	.dataa(\mem[6][67]~q ),
	.datab(\mem_used[6]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[5][67]~10_combout ),
	.cout());
defparam \mem[5][67]~10 .lut_mask = 16'hB8FF;
defparam \mem[5][67]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[5][67]~11 (
	.dataa(\mem[5][67]~q ),
	.datab(\mem[5][67]~10_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem[5][67]~11_combout ),
	.cout());
defparam \mem[5][67]~11 .lut_mask = 16'hEFFE;
defparam \mem[5][67]~11 .sum_lutc_input = "datac";

dffeas \mem[5][67] (
	.clk(clk),
	.d(\mem[5][67]~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[5][67]~q ),
	.prn(vcc));
defparam \mem[5][67] .is_wysiwyg = "true";
defparam \mem[5][67] .power_up = "low";

cycloneive_lcell_comb \mem[4][67]~8 (
	.dataa(\mem[5][67]~q ),
	.datab(\mem_used[5]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[4][67]~8_combout ),
	.cout());
defparam \mem[4][67]~8 .lut_mask = 16'hB8FF;
defparam \mem[4][67]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[4][67]~9 (
	.dataa(\mem[4][67]~q ),
	.datab(\mem[4][67]~8_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem[4][67]~9_combout ),
	.cout());
defparam \mem[4][67]~9 .lut_mask = 16'hEFFE;
defparam \mem[4][67]~9 .sum_lutc_input = "datac";

dffeas \mem[4][67] (
	.clk(clk),
	.d(\mem[4][67]~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[4][67]~q ),
	.prn(vcc));
defparam \mem[4][67] .is_wysiwyg = "true";
defparam \mem[4][67] .power_up = "low";

cycloneive_lcell_comb \mem[3][67]~6 (
	.dataa(\mem[4][67]~q ),
	.datab(\mem_used[4]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[3][67]~6_combout ),
	.cout());
defparam \mem[3][67]~6 .lut_mask = 16'hB8FF;
defparam \mem[3][67]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[3][67]~7 (
	.dataa(\mem[3][67]~q ),
	.datab(\mem[3][67]~6_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem[3][67]~7_combout ),
	.cout());
defparam \mem[3][67]~7 .lut_mask = 16'hEFFE;
defparam \mem[3][67]~7 .sum_lutc_input = "datac";

dffeas \mem[3][67] (
	.clk(clk),
	.d(\mem[3][67]~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[3][67]~q ),
	.prn(vcc));
defparam \mem[3][67] .is_wysiwyg = "true";
defparam \mem[3][67] .power_up = "low";

cycloneive_lcell_comb \mem[2][67]~4 (
	.dataa(\mem[3][67]~q ),
	.datab(\mem_used[3]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[2][67]~4_combout ),
	.cout());
defparam \mem[2][67]~4 .lut_mask = 16'hB8FF;
defparam \mem[2][67]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[2][67]~5 (
	.dataa(\mem[2][67]~q ),
	.datab(\mem[2][67]~4_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem[2][67]~5_combout ),
	.cout());
defparam \mem[2][67]~5 .lut_mask = 16'hEFFE;
defparam \mem[2][67]~5 .sum_lutc_input = "datac";

dffeas \mem[2][67] (
	.clk(clk),
	.d(\mem[2][67]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[2][67]~q ),
	.prn(vcc));
defparam \mem[2][67] .is_wysiwyg = "true";
defparam \mem[2][67] .power_up = "low";

cycloneive_lcell_comb \mem[1][67]~2 (
	.dataa(\mem[2][67]~q ),
	.datab(\mem_used[2]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[1][67]~2_combout ),
	.cout());
defparam \mem[1][67]~2 .lut_mask = 16'hB8FF;
defparam \mem[1][67]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[1][67]~3 (
	.dataa(\mem[1][67]~q ),
	.datab(\mem[1][67]~2_combout ),
	.datac(\read~0_combout ),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem[1][67]~3_combout ),
	.cout());
defparam \mem[1][67]~3 .lut_mask = 16'hEFFE;
defparam \mem[1][67]~3 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem[1][67]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem[0][67]~0 (
	.dataa(\mem[1][67]~q ),
	.datab(\mem_used[1]~q ),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem[0][67]~0_combout ),
	.cout());
defparam \mem[0][67]~0 .lut_mask = 16'hB8FF;
defparam \mem[0][67]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem[0][67]~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(out_valid),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[128]~0 (
	.dataa(\mem_used[127]~q ),
	.datab(mem_used_128),
	.datac(\read~0_combout ),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used[128]~0_combout ),
	.cout());
defparam \mem_used[128]~0 .lut_mask = 16'hEFFE;
defparam \mem_used[128]~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_2 (
	reset,
	d_write,
	write_accepted,
	sink_in_reset,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	uav_write,
	saved_grant_0,
	mem_used_1,
	uav_read,
	uav_read1,
	saved_grant_1,
	WideOr1,
	mem,
	mem1,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	write_accepted;
input 	sink_in_reset;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	uav_write;
input 	saved_grant_0;
output 	mem_used_1;
input 	uav_read;
input 	uav_read1;
input 	saved_grant_1;
input 	WideOr1;
output 	mem;
output 	mem1;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~3_combout ;
wire \mem[1][67]~q ;
wire \mem~4_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(write_accepted),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hEFFF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~1 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(mem1),
	.cout());
defparam \mem~1 .lut_mask = 16'hFFFE;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][68]~q ),
	.datab(mem1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hFAFC;
defparam \mem~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(sink_in_reset),
	.datab(WideOr1),
	.datac(mem1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~1_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_3 (
	reset,
	d_write,
	write_accepted,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	uav_write,
	uav_read,
	uav_read1,
	saved_grant_1,
	mem,
	local_read,
	mem1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	write_accepted;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
input 	uav_write;
input 	uav_read;
input 	uav_read1;
input 	saved_grant_1;
output 	mem;
input 	local_read;
output 	mem1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;
wire \mem[1][67]~q ;
wire \mem~3_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hFFFE;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~4 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(write_accepted),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(mem1),
	.cout());
defparam \mem~4 .lut_mask = 16'hEFFF;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(local_read),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hEFFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][68]~q ),
	.datab(mem),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFAFC;
defparam \mem~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(local_read),
	.datac(\mem_used[1]~0_combout ),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_4 (
	reset,
	d_write,
	write_accepted,
	read_latency_shift_reg_0,
	mem_67_0,
	uav_read,
	mem_used_1,
	av_waitrequest,
	Equal9,
	sink_ready,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	write_accepted;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	uav_read;
output 	mem_used_1;
input 	av_waitrequest;
input 	Equal9;
input 	sink_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem[1][67]~q ;
wire \mem~2_combout ;
wire \mem[0][67]~3_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~3_combout ;


dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~0_combout ),
	.cout());
defparam \mem_used[0]~0 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~1 (
	.dataa(\mem_used[0]~0_combout ),
	.datab(uav_read),
	.datac(av_waitrequest),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[0]~1_combout ),
	.cout());
defparam \mem_used[0]~1 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~1 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hB8FF;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(read_latency_shift_reg_0),
	.datac(mem_67_0),
	.datad(\mem~2_combout ),
	.cin(gnd),
	.combout(\mem[0][67]~3_combout ),
	.cout());
defparam \mem[0][67]~3 .lut_mask = 16'hFFF6;
defparam \mem[0][67]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(Equal9),
	.datac(av_waitrequest),
	.datad(uav_read),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hFFFD;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(\mem_used[1]~2_combout ),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[1]~3_combout ),
	.cout());
defparam \mem_used[1]~3 .lut_mask = 16'hDF8F;
defparam \mem_used[1]~3 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_5 (
	reset,
	mem_used_1,
	d_write,
	write_accepted,
	read_latency_shift_reg,
	read_latency_shift_reg1,
	read_latency_shift_reg_0,
	mem_67_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_used_1;
input 	d_write;
input 	write_accepted;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg1;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][67]~q ;
wire \mem~0_combout ;
wire \mem[0][67]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~2_combout ),
	.datab(read_latency_shift_reg),
	.datac(read_latency_shift_reg1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hF6F6;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(read_latency_shift_reg),
	.datab(read_latency_shift_reg1),
	.datac(mem_used_1),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hB8FF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_6 (
	d_write,
	write_accepted,
	reset,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_67_0,
	waitrequest_reset_override,
	uav_read,
	wait_latency_counter_0,
	Equal5,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	reset;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	waitrequest_reset_override;
input 	uav_read;
input 	wait_latency_counter_0;
input 	Equal5;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][67]~q ;
wire \mem~0_combout ;
wire \mem[0][67]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(uav_read),
	.datab(waitrequest_reset_override),
	.datac(Equal5),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hB8FF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_7 (
	d_write,
	write_accepted,
	reset,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_67_0,
	waitrequest_reset_override,
	uav_read,
	wait_latency_counter_1,
	Equal3,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	reset;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	waitrequest_reset_override;
input 	uav_read;
input 	wait_latency_counter_1;
input 	Equal3;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][67]~q ;
wire \mem~0_combout ;
wire \mem[0][67]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(uav_read),
	.datab(waitrequest_reset_override),
	.datac(Equal3),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hB8FF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_8 (
	clk,
	reset,
	mem_used_0,
	mem_107_0,
	out_valid1,
	WideOr0,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_22,
	out_payload_23,
	out_payload_24,
	out_payload_25,
	out_payload_26,
	out_payload_11,
	out_payload_13,
	out_payload_16,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_10,
	out_payload_9,
	out_payload_8,
	out_payload_7,
	out_payload_6,
	out_payload_20,
	out_payload_18,
	out_payload_19,
	out_payload_17,
	out_payload_21,
	out_payload_27,
	out_payload_28,
	out_payload_31,
	out_payload_30,
	out_payload_29,
	za_valid,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_22,
	za_data_23,
	za_data_24,
	za_data_25,
	za_data_26,
	za_data_11,
	za_data_13,
	za_data_16,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_10,
	za_data_9,
	za_data_8,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_18,
	za_data_19,
	za_data_17,
	za_data_21,
	za_data_27,
	za_data_28,
	za_data_31,
	za_data_30,
	za_data_29)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	mem_used_0;
input 	mem_107_0;
output 	out_valid1;
input 	WideOr0;
output 	out_payload_0;
output 	out_payload_1;
output 	out_payload_2;
output 	out_payload_3;
output 	out_payload_4;
output 	out_payload_22;
output 	out_payload_23;
output 	out_payload_24;
output 	out_payload_25;
output 	out_payload_26;
output 	out_payload_11;
output 	out_payload_13;
output 	out_payload_16;
output 	out_payload_12;
output 	out_payload_5;
output 	out_payload_14;
output 	out_payload_15;
output 	out_payload_10;
output 	out_payload_9;
output 	out_payload_8;
output 	out_payload_7;
output 	out_payload_6;
output 	out_payload_20;
output 	out_payload_18;
output 	out_payload_19;
output 	out_payload_17;
output 	out_payload_21;
output 	out_payload_27;
output 	out_payload_28;
output 	out_payload_31;
output 	out_payload_30;
output 	out_payload_29;
input 	za_valid;
input 	za_data_0;
input 	za_data_1;
input 	za_data_2;
input 	za_data_3;
input 	za_data_4;
input 	za_data_22;
input 	za_data_23;
input 	za_data_24;
input 	za_data_25;
input 	za_data_26;
input 	za_data_11;
input 	za_data_13;
input 	za_data_16;
input 	za_data_12;
input 	za_data_5;
input 	za_data_14;
input 	za_data_15;
input 	za_data_10;
input 	za_data_9;
input 	za_data_8;
input 	za_data_7;
input 	za_data_6;
input 	za_data_20;
input 	za_data_18;
input 	za_data_19;
input 	za_data_17;
input 	za_data_21;
input 	za_data_27;
input 	za_data_28;
input 	za_data_31;
input 	za_data_30;
input 	za_data_29;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \internal_out_ready~0_combout ;
wire \mem_rd_ptr[0]~1_combout ;
wire \rd_ptr[0]~q ;
wire \mem_rd_ptr[1]~0_combout ;
wire \rd_ptr[1]~q ;
wire \wr_ptr[0]~0_combout ;
wire \next_full~0_combout ;
wire \read~0_combout ;
wire \mem_rd_ptr[2]~2_combout ;
wire \rd_ptr[2]~q ;
wire \wr_ptr[2]~q ;
wire \Add0~1_combout ;
wire \next_full~1_combout ;
wire \next_full~2_combout ;
wire \full~q ;
wire \write~combout ;
wire \wr_ptr[0]~q ;
wire \Add0~0_combout ;
wire \wr_ptr[1]~q ;
wire \internal_out_valid~0_combout ;
wire \Equal0~0_combout ;
wire \internal_out_valid~1_combout ;
wire \next_empty~0_combout ;
wire \empty~q ;
wire \internal_out_valid~2_combout ;
wire \internal_out_valid~q ;
wire \mem~416_combout ;
wire \mem~160_q ;
wire \mem~417_combout ;
wire \mem~192_q ;
wire \mem~418_combout ;
wire \mem~128_q ;
wire \mem~256_combout ;
wire \mem~419_combout ;
wire \mem~224_q ;
wire \mem~257_combout ;
wire \mem~420_combout ;
wire \mem~64_q ;
wire \mem~421_combout ;
wire \mem~32_q ;
wire \mem~422_combout ;
wire \mem~0_q ;
wire \mem~258_combout ;
wire \mem~423_combout ;
wire \mem~96_q ;
wire \mem~259_combout ;
wire \mem~260_combout ;
wire \internal_out_payload[0]~q ;
wire \mem~161_q ;
wire \mem~193_q ;
wire \mem~129_q ;
wire \mem~261_combout ;
wire \mem~225_q ;
wire \mem~262_combout ;
wire \mem~65_q ;
wire \mem~33_q ;
wire \mem~1_q ;
wire \mem~263_combout ;
wire \mem~97_q ;
wire \mem~264_combout ;
wire \mem~265_combout ;
wire \internal_out_payload[1]~q ;
wire \mem~162_q ;
wire \mem~194_q ;
wire \mem~130_q ;
wire \mem~266_combout ;
wire \mem~226_q ;
wire \mem~267_combout ;
wire \mem~66_q ;
wire \mem~34_q ;
wire \mem~2_q ;
wire \mem~268_combout ;
wire \mem~98_q ;
wire \mem~269_combout ;
wire \mem~270_combout ;
wire \internal_out_payload[2]~q ;
wire \mem~163_q ;
wire \mem~195_q ;
wire \mem~131_q ;
wire \mem~271_combout ;
wire \mem~227_q ;
wire \mem~272_combout ;
wire \mem~67_q ;
wire \mem~35_q ;
wire \mem~3_q ;
wire \mem~273_combout ;
wire \mem~99_q ;
wire \mem~274_combout ;
wire \mem~275_combout ;
wire \internal_out_payload[3]~q ;
wire \mem~164_q ;
wire \mem~196_q ;
wire \mem~132_q ;
wire \mem~276_combout ;
wire \mem~228_q ;
wire \mem~277_combout ;
wire \mem~68_q ;
wire \mem~36_q ;
wire \mem~4_q ;
wire \mem~278_combout ;
wire \mem~100_q ;
wire \mem~279_combout ;
wire \mem~280_combout ;
wire \internal_out_payload[4]~q ;
wire \mem~182_q ;
wire \mem~214_q ;
wire \mem~150_q ;
wire \mem~281_combout ;
wire \mem~246_q ;
wire \mem~282_combout ;
wire \mem~86_q ;
wire \mem~54_q ;
wire \mem~22_q ;
wire \mem~283_combout ;
wire \mem~118_q ;
wire \mem~284_combout ;
wire \mem~285_combout ;
wire \internal_out_payload[22]~q ;
wire \mem~183_q ;
wire \mem~215_q ;
wire \mem~151_q ;
wire \mem~286_combout ;
wire \mem~247_q ;
wire \mem~287_combout ;
wire \mem~87_q ;
wire \mem~55_q ;
wire \mem~23_q ;
wire \mem~288_combout ;
wire \mem~119_q ;
wire \mem~289_combout ;
wire \mem~290_combout ;
wire \internal_out_payload[23]~q ;
wire \mem~184_q ;
wire \mem~216_q ;
wire \mem~152_q ;
wire \mem~291_combout ;
wire \mem~248_q ;
wire \mem~292_combout ;
wire \mem~88_q ;
wire \mem~56_q ;
wire \mem~24_q ;
wire \mem~293_combout ;
wire \mem~120_q ;
wire \mem~294_combout ;
wire \mem~295_combout ;
wire \internal_out_payload[24]~q ;
wire \mem~185_q ;
wire \mem~217_q ;
wire \mem~153_q ;
wire \mem~296_combout ;
wire \mem~249_q ;
wire \mem~297_combout ;
wire \mem~89_q ;
wire \mem~57_q ;
wire \mem~25_q ;
wire \mem~298_combout ;
wire \mem~121_q ;
wire \mem~299_combout ;
wire \mem~300_combout ;
wire \internal_out_payload[25]~q ;
wire \mem~186_q ;
wire \mem~218_q ;
wire \mem~154_q ;
wire \mem~301_combout ;
wire \mem~250_q ;
wire \mem~302_combout ;
wire \mem~90_q ;
wire \mem~58_q ;
wire \mem~26_q ;
wire \mem~303_combout ;
wire \mem~122_q ;
wire \mem~304_combout ;
wire \mem~305_combout ;
wire \internal_out_payload[26]~q ;
wire \mem~171_q ;
wire \mem~203_q ;
wire \mem~139_q ;
wire \mem~306_combout ;
wire \mem~235_q ;
wire \mem~307_combout ;
wire \mem~75_q ;
wire \mem~43_q ;
wire \mem~11_q ;
wire \mem~308_combout ;
wire \mem~107_q ;
wire \mem~309_combout ;
wire \mem~310_combout ;
wire \internal_out_payload[11]~q ;
wire \mem~173_q ;
wire \mem~205_q ;
wire \mem~141_q ;
wire \mem~311_combout ;
wire \mem~237_q ;
wire \mem~312_combout ;
wire \mem~77_q ;
wire \mem~45_q ;
wire \mem~13_q ;
wire \mem~313_combout ;
wire \mem~109_q ;
wire \mem~314_combout ;
wire \mem~315_combout ;
wire \internal_out_payload[13]~q ;
wire \mem~176_q ;
wire \mem~208_q ;
wire \mem~144_q ;
wire \mem~316_combout ;
wire \mem~240_q ;
wire \mem~317_combout ;
wire \mem~80_q ;
wire \mem~48_q ;
wire \mem~16_q ;
wire \mem~318_combout ;
wire \mem~112_q ;
wire \mem~319_combout ;
wire \mem~320_combout ;
wire \internal_out_payload[16]~q ;
wire \mem~172_q ;
wire \mem~204_q ;
wire \mem~140_q ;
wire \mem~321_combout ;
wire \mem~236_q ;
wire \mem~322_combout ;
wire \mem~76_q ;
wire \mem~44_q ;
wire \mem~12_q ;
wire \mem~323_combout ;
wire \mem~108_q ;
wire \mem~324_combout ;
wire \mem~325_combout ;
wire \internal_out_payload[12]~q ;
wire \mem~165_q ;
wire \mem~197_q ;
wire \mem~133_q ;
wire \mem~326_combout ;
wire \mem~229_q ;
wire \mem~327_combout ;
wire \mem~69_q ;
wire \mem~37_q ;
wire \mem~5_q ;
wire \mem~328_combout ;
wire \mem~101_q ;
wire \mem~329_combout ;
wire \mem~330_combout ;
wire \internal_out_payload[5]~q ;
wire \mem~174_q ;
wire \mem~206_q ;
wire \mem~142_q ;
wire \mem~331_combout ;
wire \mem~238_q ;
wire \mem~332_combout ;
wire \mem~78_q ;
wire \mem~46_q ;
wire \mem~14_q ;
wire \mem~333_combout ;
wire \mem~110_q ;
wire \mem~334_combout ;
wire \mem~335_combout ;
wire \internal_out_payload[14]~q ;
wire \mem~175_q ;
wire \mem~207_q ;
wire \mem~143_q ;
wire \mem~336_combout ;
wire \mem~239_q ;
wire \mem~337_combout ;
wire \mem~79_q ;
wire \mem~47_q ;
wire \mem~15_q ;
wire \mem~338_combout ;
wire \mem~111_q ;
wire \mem~339_combout ;
wire \mem~340_combout ;
wire \internal_out_payload[15]~q ;
wire \mem~170_q ;
wire \mem~202_q ;
wire \mem~138_q ;
wire \mem~341_combout ;
wire \mem~234_q ;
wire \mem~342_combout ;
wire \mem~74_q ;
wire \mem~42_q ;
wire \mem~10_q ;
wire \mem~343_combout ;
wire \mem~106_q ;
wire \mem~344_combout ;
wire \mem~345_combout ;
wire \internal_out_payload[10]~q ;
wire \mem~169_q ;
wire \mem~201_q ;
wire \mem~137_q ;
wire \mem~346_combout ;
wire \mem~233_q ;
wire \mem~347_combout ;
wire \mem~73_q ;
wire \mem~41_q ;
wire \mem~9_q ;
wire \mem~348_combout ;
wire \mem~105_q ;
wire \mem~349_combout ;
wire \mem~350_combout ;
wire \internal_out_payload[9]~q ;
wire \mem~168_q ;
wire \mem~200_q ;
wire \mem~136_q ;
wire \mem~351_combout ;
wire \mem~232_q ;
wire \mem~352_combout ;
wire \mem~72_q ;
wire \mem~40_q ;
wire \mem~8_q ;
wire \mem~353_combout ;
wire \mem~104_q ;
wire \mem~354_combout ;
wire \mem~355_combout ;
wire \internal_out_payload[8]~q ;
wire \mem~167_q ;
wire \mem~199_q ;
wire \mem~135_q ;
wire \mem~356_combout ;
wire \mem~231_q ;
wire \mem~357_combout ;
wire \mem~71_q ;
wire \mem~39_q ;
wire \mem~7_q ;
wire \mem~358_combout ;
wire \mem~103_q ;
wire \mem~359_combout ;
wire \mem~360_combout ;
wire \internal_out_payload[7]~q ;
wire \mem~166_q ;
wire \mem~198_q ;
wire \mem~134_q ;
wire \mem~361_combout ;
wire \mem~230_q ;
wire \mem~362_combout ;
wire \mem~70_q ;
wire \mem~38_q ;
wire \mem~6_q ;
wire \mem~363_combout ;
wire \mem~102_q ;
wire \mem~364_combout ;
wire \mem~365_combout ;
wire \internal_out_payload[6]~q ;
wire \mem~180_q ;
wire \mem~212_q ;
wire \mem~148_q ;
wire \mem~366_combout ;
wire \mem~244_q ;
wire \mem~367_combout ;
wire \mem~84_q ;
wire \mem~52_q ;
wire \mem~20_q ;
wire \mem~368_combout ;
wire \mem~116_q ;
wire \mem~369_combout ;
wire \mem~370_combout ;
wire \internal_out_payload[20]~q ;
wire \mem~178_q ;
wire \mem~210_q ;
wire \mem~146_q ;
wire \mem~371_combout ;
wire \mem~242_q ;
wire \mem~372_combout ;
wire \mem~82_q ;
wire \mem~50_q ;
wire \mem~18_q ;
wire \mem~373_combout ;
wire \mem~114_q ;
wire \mem~374_combout ;
wire \mem~375_combout ;
wire \internal_out_payload[18]~q ;
wire \mem~179_q ;
wire \mem~211_q ;
wire \mem~147_q ;
wire \mem~376_combout ;
wire \mem~243_q ;
wire \mem~377_combout ;
wire \mem~83_q ;
wire \mem~51_q ;
wire \mem~19_q ;
wire \mem~378_combout ;
wire \mem~115_q ;
wire \mem~379_combout ;
wire \mem~380_combout ;
wire \internal_out_payload[19]~q ;
wire \mem~177_q ;
wire \mem~209_q ;
wire \mem~145_q ;
wire \mem~381_combout ;
wire \mem~241_q ;
wire \mem~382_combout ;
wire \mem~81_q ;
wire \mem~49_q ;
wire \mem~17_q ;
wire \mem~383_combout ;
wire \mem~113_q ;
wire \mem~384_combout ;
wire \mem~385_combout ;
wire \internal_out_payload[17]~q ;
wire \mem~181_q ;
wire \mem~213_q ;
wire \mem~149_q ;
wire \mem~386_combout ;
wire \mem~245_q ;
wire \mem~387_combout ;
wire \mem~85_q ;
wire \mem~53_q ;
wire \mem~21_q ;
wire \mem~388_combout ;
wire \mem~117_q ;
wire \mem~389_combout ;
wire \mem~390_combout ;
wire \internal_out_payload[21]~q ;
wire \mem~187_q ;
wire \mem~219_q ;
wire \mem~155_q ;
wire \mem~391_combout ;
wire \mem~251_q ;
wire \mem~392_combout ;
wire \mem~91_q ;
wire \mem~59_q ;
wire \mem~27_q ;
wire \mem~393_combout ;
wire \mem~123_q ;
wire \mem~394_combout ;
wire \mem~395_combout ;
wire \internal_out_payload[27]~q ;
wire \mem~188_q ;
wire \mem~220_q ;
wire \mem~156_q ;
wire \mem~396_combout ;
wire \mem~252_q ;
wire \mem~397_combout ;
wire \mem~92_q ;
wire \mem~60_q ;
wire \mem~28_q ;
wire \mem~398_combout ;
wire \mem~124_q ;
wire \mem~399_combout ;
wire \mem~400_combout ;
wire \internal_out_payload[28]~q ;
wire \mem~191_q ;
wire \mem~223_q ;
wire \mem~159_q ;
wire \mem~401_combout ;
wire \mem~255_q ;
wire \mem~402_combout ;
wire \mem~95_q ;
wire \mem~63_q ;
wire \mem~31_q ;
wire \mem~403_combout ;
wire \mem~127_q ;
wire \mem~404_combout ;
wire \mem~405_combout ;
wire \internal_out_payload[31]~q ;
wire \mem~190_q ;
wire \mem~222_q ;
wire \mem~158_q ;
wire \mem~406_combout ;
wire \mem~254_q ;
wire \mem~407_combout ;
wire \mem~94_q ;
wire \mem~62_q ;
wire \mem~30_q ;
wire \mem~408_combout ;
wire \mem~126_q ;
wire \mem~409_combout ;
wire \mem~410_combout ;
wire \internal_out_payload[30]~q ;
wire \mem~189_q ;
wire \mem~221_q ;
wire \mem~157_q ;
wire \mem~411_combout ;
wire \mem~253_q ;
wire \mem~412_combout ;
wire \mem~93_q ;
wire \mem~61_q ;
wire \mem~29_q ;
wire \mem~413_combout ;
wire \mem~125_q ;
wire \mem~414_combout ;
wire \mem~415_combout ;
wire \internal_out_payload[29]~q ;


dffeas out_valid(
	.clk(clk),
	.d(\internal_out_valid~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[0] (
	.clk(clk),
	.d(\internal_out_payload[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk),
	.d(\internal_out_payload[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk),
	.d(\internal_out_payload[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas \out_payload[3] (
	.clk(clk),
	.d(\internal_out_payload[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_3),
	.prn(vcc));
defparam \out_payload[3] .is_wysiwyg = "true";
defparam \out_payload[3] .power_up = "low";

dffeas \out_payload[4] (
	.clk(clk),
	.d(\internal_out_payload[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_4),
	.prn(vcc));
defparam \out_payload[4] .is_wysiwyg = "true";
defparam \out_payload[4] .power_up = "low";

dffeas \out_payload[22] (
	.clk(clk),
	.d(\internal_out_payload[22]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_22),
	.prn(vcc));
defparam \out_payload[22] .is_wysiwyg = "true";
defparam \out_payload[22] .power_up = "low";

dffeas \out_payload[23] (
	.clk(clk),
	.d(\internal_out_payload[23]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_23),
	.prn(vcc));
defparam \out_payload[23] .is_wysiwyg = "true";
defparam \out_payload[23] .power_up = "low";

dffeas \out_payload[24] (
	.clk(clk),
	.d(\internal_out_payload[24]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_24),
	.prn(vcc));
defparam \out_payload[24] .is_wysiwyg = "true";
defparam \out_payload[24] .power_up = "low";

dffeas \out_payload[25] (
	.clk(clk),
	.d(\internal_out_payload[25]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_25),
	.prn(vcc));
defparam \out_payload[25] .is_wysiwyg = "true";
defparam \out_payload[25] .power_up = "low";

dffeas \out_payload[26] (
	.clk(clk),
	.d(\internal_out_payload[26]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_26),
	.prn(vcc));
defparam \out_payload[26] .is_wysiwyg = "true";
defparam \out_payload[26] .power_up = "low";

dffeas \out_payload[11] (
	.clk(clk),
	.d(\internal_out_payload[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_11),
	.prn(vcc));
defparam \out_payload[11] .is_wysiwyg = "true";
defparam \out_payload[11] .power_up = "low";

dffeas \out_payload[13] (
	.clk(clk),
	.d(\internal_out_payload[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_13),
	.prn(vcc));
defparam \out_payload[13] .is_wysiwyg = "true";
defparam \out_payload[13] .power_up = "low";

dffeas \out_payload[16] (
	.clk(clk),
	.d(\internal_out_payload[16]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_16),
	.prn(vcc));
defparam \out_payload[16] .is_wysiwyg = "true";
defparam \out_payload[16] .power_up = "low";

dffeas \out_payload[12] (
	.clk(clk),
	.d(\internal_out_payload[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[5] (
	.clk(clk),
	.d(\internal_out_payload[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[14] (
	.clk(clk),
	.d(\internal_out_payload[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_14),
	.prn(vcc));
defparam \out_payload[14] .is_wysiwyg = "true";
defparam \out_payload[14] .power_up = "low";

dffeas \out_payload[15] (
	.clk(clk),
	.d(\internal_out_payload[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_15),
	.prn(vcc));
defparam \out_payload[15] .is_wysiwyg = "true";
defparam \out_payload[15] .power_up = "low";

dffeas \out_payload[10] (
	.clk(clk),
	.d(\internal_out_payload[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_10),
	.prn(vcc));
defparam \out_payload[10] .is_wysiwyg = "true";
defparam \out_payload[10] .power_up = "low";

dffeas \out_payload[9] (
	.clk(clk),
	.d(\internal_out_payload[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_9),
	.prn(vcc));
defparam \out_payload[9] .is_wysiwyg = "true";
defparam \out_payload[9] .power_up = "low";

dffeas \out_payload[8] (
	.clk(clk),
	.d(\internal_out_payload[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

dffeas \out_payload[7] (
	.clk(clk),
	.d(\internal_out_payload[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[6] (
	.clk(clk),
	.d(\internal_out_payload[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

dffeas \out_payload[20] (
	.clk(clk),
	.d(\internal_out_payload[20]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_20),
	.prn(vcc));
defparam \out_payload[20] .is_wysiwyg = "true";
defparam \out_payload[20] .power_up = "low";

dffeas \out_payload[18] (
	.clk(clk),
	.d(\internal_out_payload[18]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_18),
	.prn(vcc));
defparam \out_payload[18] .is_wysiwyg = "true";
defparam \out_payload[18] .power_up = "low";

dffeas \out_payload[19] (
	.clk(clk),
	.d(\internal_out_payload[19]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_19),
	.prn(vcc));
defparam \out_payload[19] .is_wysiwyg = "true";
defparam \out_payload[19] .power_up = "low";

dffeas \out_payload[17] (
	.clk(clk),
	.d(\internal_out_payload[17]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_17),
	.prn(vcc));
defparam \out_payload[17] .is_wysiwyg = "true";
defparam \out_payload[17] .power_up = "low";

dffeas \out_payload[21] (
	.clk(clk),
	.d(\internal_out_payload[21]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_21),
	.prn(vcc));
defparam \out_payload[21] .is_wysiwyg = "true";
defparam \out_payload[21] .power_up = "low";

dffeas \out_payload[27] (
	.clk(clk),
	.d(\internal_out_payload[27]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_27),
	.prn(vcc));
defparam \out_payload[27] .is_wysiwyg = "true";
defparam \out_payload[27] .power_up = "low";

dffeas \out_payload[28] (
	.clk(clk),
	.d(\internal_out_payload[28]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_28),
	.prn(vcc));
defparam \out_payload[28] .is_wysiwyg = "true";
defparam \out_payload[28] .power_up = "low";

dffeas \out_payload[31] (
	.clk(clk),
	.d(\internal_out_payload[31]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_31),
	.prn(vcc));
defparam \out_payload[31] .is_wysiwyg = "true";
defparam \out_payload[31] .power_up = "low";

dffeas \out_payload[30] (
	.clk(clk),
	.d(\internal_out_payload[30]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_30),
	.prn(vcc));
defparam \out_payload[30] .is_wysiwyg = "true";
defparam \out_payload[30] .power_up = "low";

dffeas \out_payload[29] (
	.clk(clk),
	.d(\internal_out_payload[29]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_29),
	.prn(vcc));
defparam \out_payload[29] .is_wysiwyg = "true";
defparam \out_payload[29] .power_up = "low";

cycloneive_lcell_comb \internal_out_ready~0 (
	.dataa(mem_used_0),
	.datab(mem_107_0),
	.datac(WideOr0),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_ready~0_combout ),
	.cout());
defparam \internal_out_ready~0 .lut_mask = 16'h7FFF;
defparam \internal_out_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[0]~1 (
	.dataa(gnd),
	.datab(\rd_ptr[0]~q ),
	.datac(\internal_out_valid~q ),
	.datad(\internal_out_ready~0_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[0]~1_combout ),
	.cout());
defparam \mem_rd_ptr[0]~1 .lut_mask = 16'hC33C;
defparam \mem_rd_ptr[0]~1 .sum_lutc_input = "datac";

dffeas \rd_ptr[0] (
	.clk(clk),
	.d(\mem_rd_ptr[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[0]~q ),
	.prn(vcc));
defparam \rd_ptr[0] .is_wysiwyg = "true";
defparam \rd_ptr[0] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[1]~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\internal_out_valid~q ),
	.datac(\internal_out_ready~0_combout ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[1]~0_combout ),
	.cout());
defparam \mem_rd_ptr[1]~0 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[1]~0 .sum_lutc_input = "datac";

dffeas \rd_ptr[1] (
	.clk(clk),
	.d(\mem_rd_ptr[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[1]~q ),
	.prn(vcc));
defparam \rd_ptr[1] .is_wysiwyg = "true";
defparam \rd_ptr[1] .power_up = "low";

cycloneive_lcell_comb \wr_ptr[0]~0 (
	.dataa(\wr_ptr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_ptr[0]~0_combout ),
	.cout());
defparam \wr_ptr[0]~0 .lut_mask = 16'h5555;
defparam \wr_ptr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\next_full~0_combout ),
	.cout());
defparam \next_full~0 .lut_mask = 16'h6996;
defparam \next_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(\internal_out_valid~q ),
	.datab(\internal_out_ready~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hEEEE;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[2]~2 (
	.dataa(\rd_ptr[2]~q ),
	.datab(\read~0_combout ),
	.datac(\rd_ptr[1]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[2]~2_combout ),
	.cout());
defparam \mem_rd_ptr[2]~2 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[2]~2 .sum_lutc_input = "datac";

dffeas \rd_ptr[2] (
	.clk(clk),
	.d(\mem_rd_ptr[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[2]~q ),
	.prn(vcc));
defparam \rd_ptr[2] .is_wysiwyg = "true";
defparam \rd_ptr[2] .power_up = "low";

dffeas \wr_ptr[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_ptr[2] .is_wysiwyg = "true";
defparam \wr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'hC33C;
defparam \Add0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~1 (
	.dataa(za_valid),
	.datab(\next_full~0_combout ),
	.datac(\rd_ptr[2]~q ),
	.datad(\Add0~1_combout ),
	.cin(gnd),
	.combout(\next_full~1_combout ),
	.cout());
defparam \next_full~1 .lut_mask = 16'hEFFE;
defparam \next_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~2 (
	.dataa(\full~q ),
	.datab(\next_full~1_combout ),
	.datac(\internal_out_valid~q ),
	.datad(\internal_out_ready~0_combout ),
	.cin(gnd),
	.combout(\next_full~2_combout ),
	.cout());
defparam \next_full~2 .lut_mask = 16'hEFFF;
defparam \next_full~2 .sum_lutc_input = "datac";

dffeas full(
	.clk(clk),
	.d(\next_full~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\full~q ),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

cycloneive_lcell_comb write(
	.dataa(za_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(\full~q ),
	.cin(gnd),
	.combout(\write~combout ),
	.cout());
defparam write.lut_mask = 16'hAAFF;
defparam write.sum_lutc_input = "datac";

dffeas \wr_ptr[0] (
	.clk(clk),
	.d(\wr_ptr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_ptr[0] .is_wysiwyg = "true";
defparam \wr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \wr_ptr[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_ptr[1] .is_wysiwyg = "true";
defparam \wr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \internal_out_valid~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\internal_out_valid~0_combout ),
	.cout());
defparam \internal_out_valid~0 .lut_mask = 16'h6996;
defparam \internal_out_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\rd_ptr[0]~q ),
	.datac(\wr_ptr[2]~q ),
	.datad(\rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_valid~1 (
	.dataa(\internal_out_valid~q ),
	.datab(\internal_out_ready~0_combout ),
	.datac(\internal_out_valid~0_combout ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~1_combout ),
	.cout());
defparam \internal_out_valid~1 .lut_mask = 16'hFEFF;
defparam \internal_out_valid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_empty~0 (
	.dataa(\read~0_combout ),
	.datab(\internal_out_valid~1_combout ),
	.datac(\empty~q ),
	.datad(\write~combout ),
	.cin(gnd),
	.combout(\next_empty~0_combout ),
	.cout());
defparam \next_empty~0 .lut_mask = 16'hFFF7;
defparam \next_empty~0 .sum_lutc_input = "datac";

dffeas empty(
	.clk(clk),
	.d(\next_empty~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

cycloneive_lcell_comb \internal_out_valid~2 (
	.dataa(\internal_out_valid~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\empty~q ),
	.cin(gnd),
	.combout(\internal_out_valid~2_combout ),
	.cout());
defparam \internal_out_valid~2 .lut_mask = 16'hFF55;
defparam \internal_out_valid~2 .sum_lutc_input = "datac";

dffeas internal_out_valid(
	.clk(clk),
	.d(\internal_out_valid~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_valid~q ),
	.prn(vcc));
defparam internal_out_valid.is_wysiwyg = "true";
defparam internal_out_valid.power_up = "low";

cycloneive_lcell_comb \mem~416 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~416_combout ),
	.cout());
defparam \mem~416 .lut_mask = 16'hFEFF;
defparam \mem~416 .sum_lutc_input = "datac";

dffeas \mem~160 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~160_q ),
	.prn(vcc));
defparam \mem~160 .is_wysiwyg = "true";
defparam \mem~160 .power_up = "low";

cycloneive_lcell_comb \mem~417 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem~417_combout ),
	.cout());
defparam \mem~417 .lut_mask = 16'hFEFF;
defparam \mem~417 .sum_lutc_input = "datac";

dffeas \mem~192 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~192_q ),
	.prn(vcc));
defparam \mem~192 .is_wysiwyg = "true";
defparam \mem~192 .power_up = "low";

cycloneive_lcell_comb \mem~418 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~418_combout ),
	.cout());
defparam \mem~418 .lut_mask = 16'hEFFF;
defparam \mem~418 .sum_lutc_input = "datac";

dffeas \mem~128 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~128_q ),
	.prn(vcc));
defparam \mem~128 .is_wysiwyg = "true";
defparam \mem~128 .power_up = "low";

cycloneive_lcell_comb \mem~256 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~192_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~128_q ),
	.cin(gnd),
	.combout(\mem~256_combout ),
	.cout());
defparam \mem~256 .lut_mask = 16'hFFDE;
defparam \mem~256 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~419 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\write~combout ),
	.cin(gnd),
	.combout(\mem~419_combout ),
	.cout());
defparam \mem~419 .lut_mask = 16'hFFFE;
defparam \mem~419 .sum_lutc_input = "datac";

dffeas \mem~224 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~224_q ),
	.prn(vcc));
defparam \mem~224 .is_wysiwyg = "true";
defparam \mem~224 .power_up = "low";

cycloneive_lcell_comb \mem~257 (
	.dataa(\mem~160_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~256_combout ),
	.datad(\mem~224_q ),
	.cin(gnd),
	.combout(\mem~257_combout ),
	.cout());
defparam \mem~257 .lut_mask = 16'hFFBE;
defparam \mem~257 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~420 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem~420_combout ),
	.cout());
defparam \mem~420 .lut_mask = 16'hEFFF;
defparam \mem~420 .sum_lutc_input = "datac";

dffeas \mem~64 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~64_q ),
	.prn(vcc));
defparam \mem~64 .is_wysiwyg = "true";
defparam \mem~64 .power_up = "low";

cycloneive_lcell_comb \mem~421 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~421_combout ),
	.cout());
defparam \mem~421 .lut_mask = 16'hEFFF;
defparam \mem~421 .sum_lutc_input = "datac";

dffeas \mem~32 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~32_q ),
	.prn(vcc));
defparam \mem~32 .is_wysiwyg = "true";
defparam \mem~32 .power_up = "low";

cycloneive_lcell_comb \mem~422 (
	.dataa(\write~combout ),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~422_combout ),
	.cout());
defparam \mem~422 .lut_mask = 16'hBFFF;
defparam \mem~422 .sum_lutc_input = "datac";

dffeas \mem~0 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~0_q ),
	.prn(vcc));
defparam \mem~0 .is_wysiwyg = "true";
defparam \mem~0 .power_up = "low";

cycloneive_lcell_comb \mem~258 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~32_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~0_q ),
	.cin(gnd),
	.combout(\mem~258_combout ),
	.cout());
defparam \mem~258 .lut_mask = 16'hFFDE;
defparam \mem~258 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~423 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[2]~q ),
	.cin(gnd),
	.combout(\mem~423_combout ),
	.cout());
defparam \mem~423 .lut_mask = 16'hFEFF;
defparam \mem~423 .sum_lutc_input = "datac";

dffeas \mem~96 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~96_q ),
	.prn(vcc));
defparam \mem~96 .is_wysiwyg = "true";
defparam \mem~96 .power_up = "low";

cycloneive_lcell_comb \mem~259 (
	.dataa(\mem~64_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~258_combout ),
	.datad(\mem~96_q ),
	.cin(gnd),
	.combout(\mem~259_combout ),
	.cout());
defparam \mem~259 .lut_mask = 16'hFFBE;
defparam \mem~259 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~260 (
	.dataa(\mem~257_combout ),
	.datab(\mem~259_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~260_combout ),
	.cout());
defparam \mem~260 .lut_mask = 16'hAACC;
defparam \mem~260 .sum_lutc_input = "datac";

dffeas \internal_out_payload[0] (
	.clk(clk),
	.d(\mem~260_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[0]~q ),
	.prn(vcc));
defparam \internal_out_payload[0] .is_wysiwyg = "true";
defparam \internal_out_payload[0] .power_up = "low";

dffeas \mem~161 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~161_q ),
	.prn(vcc));
defparam \mem~161 .is_wysiwyg = "true";
defparam \mem~161 .power_up = "low";

dffeas \mem~193 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~193_q ),
	.prn(vcc));
defparam \mem~193 .is_wysiwyg = "true";
defparam \mem~193 .power_up = "low";

dffeas \mem~129 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~129_q ),
	.prn(vcc));
defparam \mem~129 .is_wysiwyg = "true";
defparam \mem~129 .power_up = "low";

cycloneive_lcell_comb \mem~261 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~193_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~129_q ),
	.cin(gnd),
	.combout(\mem~261_combout ),
	.cout());
defparam \mem~261 .lut_mask = 16'hFFDE;
defparam \mem~261 .sum_lutc_input = "datac";

dffeas \mem~225 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~225_q ),
	.prn(vcc));
defparam \mem~225 .is_wysiwyg = "true";
defparam \mem~225 .power_up = "low";

cycloneive_lcell_comb \mem~262 (
	.dataa(\mem~161_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~261_combout ),
	.datad(\mem~225_q ),
	.cin(gnd),
	.combout(\mem~262_combout ),
	.cout());
defparam \mem~262 .lut_mask = 16'hFFBE;
defparam \mem~262 .sum_lutc_input = "datac";

dffeas \mem~65 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~65_q ),
	.prn(vcc));
defparam \mem~65 .is_wysiwyg = "true";
defparam \mem~65 .power_up = "low";

dffeas \mem~33 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~33_q ),
	.prn(vcc));
defparam \mem~33 .is_wysiwyg = "true";
defparam \mem~33 .power_up = "low";

dffeas \mem~1 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~1_q ),
	.prn(vcc));
defparam \mem~1 .is_wysiwyg = "true";
defparam \mem~1 .power_up = "low";

cycloneive_lcell_comb \mem~263 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~33_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~1_q ),
	.cin(gnd),
	.combout(\mem~263_combout ),
	.cout());
defparam \mem~263 .lut_mask = 16'hFFDE;
defparam \mem~263 .sum_lutc_input = "datac";

dffeas \mem~97 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~97_q ),
	.prn(vcc));
defparam \mem~97 .is_wysiwyg = "true";
defparam \mem~97 .power_up = "low";

cycloneive_lcell_comb \mem~264 (
	.dataa(\mem~65_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~263_combout ),
	.datad(\mem~97_q ),
	.cin(gnd),
	.combout(\mem~264_combout ),
	.cout());
defparam \mem~264 .lut_mask = 16'hFFBE;
defparam \mem~264 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~265 (
	.dataa(\mem~262_combout ),
	.datab(\mem~264_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~265_combout ),
	.cout());
defparam \mem~265 .lut_mask = 16'hAACC;
defparam \mem~265 .sum_lutc_input = "datac";

dffeas \internal_out_payload[1] (
	.clk(clk),
	.d(\mem~265_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[1]~q ),
	.prn(vcc));
defparam \internal_out_payload[1] .is_wysiwyg = "true";
defparam \internal_out_payload[1] .power_up = "low";

dffeas \mem~162 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~162_q ),
	.prn(vcc));
defparam \mem~162 .is_wysiwyg = "true";
defparam \mem~162 .power_up = "low";

dffeas \mem~194 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~194_q ),
	.prn(vcc));
defparam \mem~194 .is_wysiwyg = "true";
defparam \mem~194 .power_up = "low";

dffeas \mem~130 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~130_q ),
	.prn(vcc));
defparam \mem~130 .is_wysiwyg = "true";
defparam \mem~130 .power_up = "low";

cycloneive_lcell_comb \mem~266 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~194_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~130_q ),
	.cin(gnd),
	.combout(\mem~266_combout ),
	.cout());
defparam \mem~266 .lut_mask = 16'hFFDE;
defparam \mem~266 .sum_lutc_input = "datac";

dffeas \mem~226 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~226_q ),
	.prn(vcc));
defparam \mem~226 .is_wysiwyg = "true";
defparam \mem~226 .power_up = "low";

cycloneive_lcell_comb \mem~267 (
	.dataa(\mem~162_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~266_combout ),
	.datad(\mem~226_q ),
	.cin(gnd),
	.combout(\mem~267_combout ),
	.cout());
defparam \mem~267 .lut_mask = 16'hFFBE;
defparam \mem~267 .sum_lutc_input = "datac";

dffeas \mem~66 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~66_q ),
	.prn(vcc));
defparam \mem~66 .is_wysiwyg = "true";
defparam \mem~66 .power_up = "low";

dffeas \mem~34 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~34_q ),
	.prn(vcc));
defparam \mem~34 .is_wysiwyg = "true";
defparam \mem~34 .power_up = "low";

dffeas \mem~2 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~2_q ),
	.prn(vcc));
defparam \mem~2 .is_wysiwyg = "true";
defparam \mem~2 .power_up = "low";

cycloneive_lcell_comb \mem~268 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~34_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~2_q ),
	.cin(gnd),
	.combout(\mem~268_combout ),
	.cout());
defparam \mem~268 .lut_mask = 16'hFFDE;
defparam \mem~268 .sum_lutc_input = "datac";

dffeas \mem~98 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~98_q ),
	.prn(vcc));
defparam \mem~98 .is_wysiwyg = "true";
defparam \mem~98 .power_up = "low";

cycloneive_lcell_comb \mem~269 (
	.dataa(\mem~66_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~268_combout ),
	.datad(\mem~98_q ),
	.cin(gnd),
	.combout(\mem~269_combout ),
	.cout());
defparam \mem~269 .lut_mask = 16'hFFBE;
defparam \mem~269 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~270 (
	.dataa(\mem~267_combout ),
	.datab(\mem~269_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~270_combout ),
	.cout());
defparam \mem~270 .lut_mask = 16'hAACC;
defparam \mem~270 .sum_lutc_input = "datac";

dffeas \internal_out_payload[2] (
	.clk(clk),
	.d(\mem~270_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[2]~q ),
	.prn(vcc));
defparam \internal_out_payload[2] .is_wysiwyg = "true";
defparam \internal_out_payload[2] .power_up = "low";

dffeas \mem~163 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~163_q ),
	.prn(vcc));
defparam \mem~163 .is_wysiwyg = "true";
defparam \mem~163 .power_up = "low";

dffeas \mem~195 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~195_q ),
	.prn(vcc));
defparam \mem~195 .is_wysiwyg = "true";
defparam \mem~195 .power_up = "low";

dffeas \mem~131 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~131_q ),
	.prn(vcc));
defparam \mem~131 .is_wysiwyg = "true";
defparam \mem~131 .power_up = "low";

cycloneive_lcell_comb \mem~271 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~195_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~131_q ),
	.cin(gnd),
	.combout(\mem~271_combout ),
	.cout());
defparam \mem~271 .lut_mask = 16'hFFDE;
defparam \mem~271 .sum_lutc_input = "datac";

dffeas \mem~227 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~227_q ),
	.prn(vcc));
defparam \mem~227 .is_wysiwyg = "true";
defparam \mem~227 .power_up = "low";

cycloneive_lcell_comb \mem~272 (
	.dataa(\mem~163_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~271_combout ),
	.datad(\mem~227_q ),
	.cin(gnd),
	.combout(\mem~272_combout ),
	.cout());
defparam \mem~272 .lut_mask = 16'hFFBE;
defparam \mem~272 .sum_lutc_input = "datac";

dffeas \mem~67 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~67_q ),
	.prn(vcc));
defparam \mem~67 .is_wysiwyg = "true";
defparam \mem~67 .power_up = "low";

dffeas \mem~35 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~35_q ),
	.prn(vcc));
defparam \mem~35 .is_wysiwyg = "true";
defparam \mem~35 .power_up = "low";

dffeas \mem~3 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~3_q ),
	.prn(vcc));
defparam \mem~3 .is_wysiwyg = "true";
defparam \mem~3 .power_up = "low";

cycloneive_lcell_comb \mem~273 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~35_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~3_q ),
	.cin(gnd),
	.combout(\mem~273_combout ),
	.cout());
defparam \mem~273 .lut_mask = 16'hFFDE;
defparam \mem~273 .sum_lutc_input = "datac";

dffeas \mem~99 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~99_q ),
	.prn(vcc));
defparam \mem~99 .is_wysiwyg = "true";
defparam \mem~99 .power_up = "low";

cycloneive_lcell_comb \mem~274 (
	.dataa(\mem~67_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~273_combout ),
	.datad(\mem~99_q ),
	.cin(gnd),
	.combout(\mem~274_combout ),
	.cout());
defparam \mem~274 .lut_mask = 16'hFFBE;
defparam \mem~274 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~275 (
	.dataa(\mem~272_combout ),
	.datab(\mem~274_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~275_combout ),
	.cout());
defparam \mem~275 .lut_mask = 16'hAACC;
defparam \mem~275 .sum_lutc_input = "datac";

dffeas \internal_out_payload[3] (
	.clk(clk),
	.d(\mem~275_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[3]~q ),
	.prn(vcc));
defparam \internal_out_payload[3] .is_wysiwyg = "true";
defparam \internal_out_payload[3] .power_up = "low";

dffeas \mem~164 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~164_q ),
	.prn(vcc));
defparam \mem~164 .is_wysiwyg = "true";
defparam \mem~164 .power_up = "low";

dffeas \mem~196 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~196_q ),
	.prn(vcc));
defparam \mem~196 .is_wysiwyg = "true";
defparam \mem~196 .power_up = "low";

dffeas \mem~132 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~132_q ),
	.prn(vcc));
defparam \mem~132 .is_wysiwyg = "true";
defparam \mem~132 .power_up = "low";

cycloneive_lcell_comb \mem~276 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~196_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~132_q ),
	.cin(gnd),
	.combout(\mem~276_combout ),
	.cout());
defparam \mem~276 .lut_mask = 16'hFFDE;
defparam \mem~276 .sum_lutc_input = "datac";

dffeas \mem~228 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~228_q ),
	.prn(vcc));
defparam \mem~228 .is_wysiwyg = "true";
defparam \mem~228 .power_up = "low";

cycloneive_lcell_comb \mem~277 (
	.dataa(\mem~164_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~276_combout ),
	.datad(\mem~228_q ),
	.cin(gnd),
	.combout(\mem~277_combout ),
	.cout());
defparam \mem~277 .lut_mask = 16'hFFBE;
defparam \mem~277 .sum_lutc_input = "datac";

dffeas \mem~68 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~68_q ),
	.prn(vcc));
defparam \mem~68 .is_wysiwyg = "true";
defparam \mem~68 .power_up = "low";

dffeas \mem~36 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~36_q ),
	.prn(vcc));
defparam \mem~36 .is_wysiwyg = "true";
defparam \mem~36 .power_up = "low";

dffeas \mem~4 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~4_q ),
	.prn(vcc));
defparam \mem~4 .is_wysiwyg = "true";
defparam \mem~4 .power_up = "low";

cycloneive_lcell_comb \mem~278 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~36_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~4_q ),
	.cin(gnd),
	.combout(\mem~278_combout ),
	.cout());
defparam \mem~278 .lut_mask = 16'hFFDE;
defparam \mem~278 .sum_lutc_input = "datac";

dffeas \mem~100 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~100_q ),
	.prn(vcc));
defparam \mem~100 .is_wysiwyg = "true";
defparam \mem~100 .power_up = "low";

cycloneive_lcell_comb \mem~279 (
	.dataa(\mem~68_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~278_combout ),
	.datad(\mem~100_q ),
	.cin(gnd),
	.combout(\mem~279_combout ),
	.cout());
defparam \mem~279 .lut_mask = 16'hFFBE;
defparam \mem~279 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~280 (
	.dataa(\mem~277_combout ),
	.datab(\mem~279_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~280_combout ),
	.cout());
defparam \mem~280 .lut_mask = 16'hAACC;
defparam \mem~280 .sum_lutc_input = "datac";

dffeas \internal_out_payload[4] (
	.clk(clk),
	.d(\mem~280_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[4]~q ),
	.prn(vcc));
defparam \internal_out_payload[4] .is_wysiwyg = "true";
defparam \internal_out_payload[4] .power_up = "low";

dffeas \mem~182 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~182_q ),
	.prn(vcc));
defparam \mem~182 .is_wysiwyg = "true";
defparam \mem~182 .power_up = "low";

dffeas \mem~214 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~214_q ),
	.prn(vcc));
defparam \mem~214 .is_wysiwyg = "true";
defparam \mem~214 .power_up = "low";

dffeas \mem~150 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~150_q ),
	.prn(vcc));
defparam \mem~150 .is_wysiwyg = "true";
defparam \mem~150 .power_up = "low";

cycloneive_lcell_comb \mem~281 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~214_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~150_q ),
	.cin(gnd),
	.combout(\mem~281_combout ),
	.cout());
defparam \mem~281 .lut_mask = 16'hFFDE;
defparam \mem~281 .sum_lutc_input = "datac";

dffeas \mem~246 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~246_q ),
	.prn(vcc));
defparam \mem~246 .is_wysiwyg = "true";
defparam \mem~246 .power_up = "low";

cycloneive_lcell_comb \mem~282 (
	.dataa(\mem~182_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~281_combout ),
	.datad(\mem~246_q ),
	.cin(gnd),
	.combout(\mem~282_combout ),
	.cout());
defparam \mem~282 .lut_mask = 16'hFFBE;
defparam \mem~282 .sum_lutc_input = "datac";

dffeas \mem~86 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~86_q ),
	.prn(vcc));
defparam \mem~86 .is_wysiwyg = "true";
defparam \mem~86 .power_up = "low";

dffeas \mem~54 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~54_q ),
	.prn(vcc));
defparam \mem~54 .is_wysiwyg = "true";
defparam \mem~54 .power_up = "low";

dffeas \mem~22 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~22_q ),
	.prn(vcc));
defparam \mem~22 .is_wysiwyg = "true";
defparam \mem~22 .power_up = "low";

cycloneive_lcell_comb \mem~283 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~54_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~22_q ),
	.cin(gnd),
	.combout(\mem~283_combout ),
	.cout());
defparam \mem~283 .lut_mask = 16'hFFDE;
defparam \mem~283 .sum_lutc_input = "datac";

dffeas \mem~118 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~118_q ),
	.prn(vcc));
defparam \mem~118 .is_wysiwyg = "true";
defparam \mem~118 .power_up = "low";

cycloneive_lcell_comb \mem~284 (
	.dataa(\mem~86_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~283_combout ),
	.datad(\mem~118_q ),
	.cin(gnd),
	.combout(\mem~284_combout ),
	.cout());
defparam \mem~284 .lut_mask = 16'hFFBE;
defparam \mem~284 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~285 (
	.dataa(\mem~282_combout ),
	.datab(\mem~284_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~285_combout ),
	.cout());
defparam \mem~285 .lut_mask = 16'hAACC;
defparam \mem~285 .sum_lutc_input = "datac";

dffeas \internal_out_payload[22] (
	.clk(clk),
	.d(\mem~285_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[22]~q ),
	.prn(vcc));
defparam \internal_out_payload[22] .is_wysiwyg = "true";
defparam \internal_out_payload[22] .power_up = "low";

dffeas \mem~183 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~183_q ),
	.prn(vcc));
defparam \mem~183 .is_wysiwyg = "true";
defparam \mem~183 .power_up = "low";

dffeas \mem~215 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~215_q ),
	.prn(vcc));
defparam \mem~215 .is_wysiwyg = "true";
defparam \mem~215 .power_up = "low";

dffeas \mem~151 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~151_q ),
	.prn(vcc));
defparam \mem~151 .is_wysiwyg = "true";
defparam \mem~151 .power_up = "low";

cycloneive_lcell_comb \mem~286 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~215_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~151_q ),
	.cin(gnd),
	.combout(\mem~286_combout ),
	.cout());
defparam \mem~286 .lut_mask = 16'hFFDE;
defparam \mem~286 .sum_lutc_input = "datac";

dffeas \mem~247 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~247_q ),
	.prn(vcc));
defparam \mem~247 .is_wysiwyg = "true";
defparam \mem~247 .power_up = "low";

cycloneive_lcell_comb \mem~287 (
	.dataa(\mem~183_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~286_combout ),
	.datad(\mem~247_q ),
	.cin(gnd),
	.combout(\mem~287_combout ),
	.cout());
defparam \mem~287 .lut_mask = 16'hFFBE;
defparam \mem~287 .sum_lutc_input = "datac";

dffeas \mem~87 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~87_q ),
	.prn(vcc));
defparam \mem~87 .is_wysiwyg = "true";
defparam \mem~87 .power_up = "low";

dffeas \mem~55 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~55_q ),
	.prn(vcc));
defparam \mem~55 .is_wysiwyg = "true";
defparam \mem~55 .power_up = "low";

dffeas \mem~23 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~23_q ),
	.prn(vcc));
defparam \mem~23 .is_wysiwyg = "true";
defparam \mem~23 .power_up = "low";

cycloneive_lcell_comb \mem~288 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~55_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~23_q ),
	.cin(gnd),
	.combout(\mem~288_combout ),
	.cout());
defparam \mem~288 .lut_mask = 16'hFFDE;
defparam \mem~288 .sum_lutc_input = "datac";

dffeas \mem~119 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~119_q ),
	.prn(vcc));
defparam \mem~119 .is_wysiwyg = "true";
defparam \mem~119 .power_up = "low";

cycloneive_lcell_comb \mem~289 (
	.dataa(\mem~87_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~288_combout ),
	.datad(\mem~119_q ),
	.cin(gnd),
	.combout(\mem~289_combout ),
	.cout());
defparam \mem~289 .lut_mask = 16'hFFBE;
defparam \mem~289 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~290 (
	.dataa(\mem~287_combout ),
	.datab(\mem~289_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~290_combout ),
	.cout());
defparam \mem~290 .lut_mask = 16'hAACC;
defparam \mem~290 .sum_lutc_input = "datac";

dffeas \internal_out_payload[23] (
	.clk(clk),
	.d(\mem~290_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[23]~q ),
	.prn(vcc));
defparam \internal_out_payload[23] .is_wysiwyg = "true";
defparam \internal_out_payload[23] .power_up = "low";

dffeas \mem~184 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~184_q ),
	.prn(vcc));
defparam \mem~184 .is_wysiwyg = "true";
defparam \mem~184 .power_up = "low";

dffeas \mem~216 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~216_q ),
	.prn(vcc));
defparam \mem~216 .is_wysiwyg = "true";
defparam \mem~216 .power_up = "low";

dffeas \mem~152 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~152_q ),
	.prn(vcc));
defparam \mem~152 .is_wysiwyg = "true";
defparam \mem~152 .power_up = "low";

cycloneive_lcell_comb \mem~291 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~216_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~152_q ),
	.cin(gnd),
	.combout(\mem~291_combout ),
	.cout());
defparam \mem~291 .lut_mask = 16'hFFDE;
defparam \mem~291 .sum_lutc_input = "datac";

dffeas \mem~248 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~248_q ),
	.prn(vcc));
defparam \mem~248 .is_wysiwyg = "true";
defparam \mem~248 .power_up = "low";

cycloneive_lcell_comb \mem~292 (
	.dataa(\mem~184_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~291_combout ),
	.datad(\mem~248_q ),
	.cin(gnd),
	.combout(\mem~292_combout ),
	.cout());
defparam \mem~292 .lut_mask = 16'hFFBE;
defparam \mem~292 .sum_lutc_input = "datac";

dffeas \mem~88 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~88_q ),
	.prn(vcc));
defparam \mem~88 .is_wysiwyg = "true";
defparam \mem~88 .power_up = "low";

dffeas \mem~56 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~56_q ),
	.prn(vcc));
defparam \mem~56 .is_wysiwyg = "true";
defparam \mem~56 .power_up = "low";

dffeas \mem~24 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~24_q ),
	.prn(vcc));
defparam \mem~24 .is_wysiwyg = "true";
defparam \mem~24 .power_up = "low";

cycloneive_lcell_comb \mem~293 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~56_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~24_q ),
	.cin(gnd),
	.combout(\mem~293_combout ),
	.cout());
defparam \mem~293 .lut_mask = 16'hFFDE;
defparam \mem~293 .sum_lutc_input = "datac";

dffeas \mem~120 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~120_q ),
	.prn(vcc));
defparam \mem~120 .is_wysiwyg = "true";
defparam \mem~120 .power_up = "low";

cycloneive_lcell_comb \mem~294 (
	.dataa(\mem~88_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~293_combout ),
	.datad(\mem~120_q ),
	.cin(gnd),
	.combout(\mem~294_combout ),
	.cout());
defparam \mem~294 .lut_mask = 16'hFFBE;
defparam \mem~294 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~295 (
	.dataa(\mem~292_combout ),
	.datab(\mem~294_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~295_combout ),
	.cout());
defparam \mem~295 .lut_mask = 16'hAACC;
defparam \mem~295 .sum_lutc_input = "datac";

dffeas \internal_out_payload[24] (
	.clk(clk),
	.d(\mem~295_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[24]~q ),
	.prn(vcc));
defparam \internal_out_payload[24] .is_wysiwyg = "true";
defparam \internal_out_payload[24] .power_up = "low";

dffeas \mem~185 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~185_q ),
	.prn(vcc));
defparam \mem~185 .is_wysiwyg = "true";
defparam \mem~185 .power_up = "low";

dffeas \mem~217 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~217_q ),
	.prn(vcc));
defparam \mem~217 .is_wysiwyg = "true";
defparam \mem~217 .power_up = "low";

dffeas \mem~153 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~153_q ),
	.prn(vcc));
defparam \mem~153 .is_wysiwyg = "true";
defparam \mem~153 .power_up = "low";

cycloneive_lcell_comb \mem~296 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~217_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~153_q ),
	.cin(gnd),
	.combout(\mem~296_combout ),
	.cout());
defparam \mem~296 .lut_mask = 16'hFFDE;
defparam \mem~296 .sum_lutc_input = "datac";

dffeas \mem~249 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~249_q ),
	.prn(vcc));
defparam \mem~249 .is_wysiwyg = "true";
defparam \mem~249 .power_up = "low";

cycloneive_lcell_comb \mem~297 (
	.dataa(\mem~185_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~296_combout ),
	.datad(\mem~249_q ),
	.cin(gnd),
	.combout(\mem~297_combout ),
	.cout());
defparam \mem~297 .lut_mask = 16'hFFBE;
defparam \mem~297 .sum_lutc_input = "datac";

dffeas \mem~89 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~89_q ),
	.prn(vcc));
defparam \mem~89 .is_wysiwyg = "true";
defparam \mem~89 .power_up = "low";

dffeas \mem~57 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~57_q ),
	.prn(vcc));
defparam \mem~57 .is_wysiwyg = "true";
defparam \mem~57 .power_up = "low";

dffeas \mem~25 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~25_q ),
	.prn(vcc));
defparam \mem~25 .is_wysiwyg = "true";
defparam \mem~25 .power_up = "low";

cycloneive_lcell_comb \mem~298 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~57_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~25_q ),
	.cin(gnd),
	.combout(\mem~298_combout ),
	.cout());
defparam \mem~298 .lut_mask = 16'hFFDE;
defparam \mem~298 .sum_lutc_input = "datac";

dffeas \mem~121 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~121_q ),
	.prn(vcc));
defparam \mem~121 .is_wysiwyg = "true";
defparam \mem~121 .power_up = "low";

cycloneive_lcell_comb \mem~299 (
	.dataa(\mem~89_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~298_combout ),
	.datad(\mem~121_q ),
	.cin(gnd),
	.combout(\mem~299_combout ),
	.cout());
defparam \mem~299 .lut_mask = 16'hFFBE;
defparam \mem~299 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~300 (
	.dataa(\mem~297_combout ),
	.datab(\mem~299_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~300_combout ),
	.cout());
defparam \mem~300 .lut_mask = 16'hAACC;
defparam \mem~300 .sum_lutc_input = "datac";

dffeas \internal_out_payload[25] (
	.clk(clk),
	.d(\mem~300_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[25]~q ),
	.prn(vcc));
defparam \internal_out_payload[25] .is_wysiwyg = "true";
defparam \internal_out_payload[25] .power_up = "low";

dffeas \mem~186 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~186_q ),
	.prn(vcc));
defparam \mem~186 .is_wysiwyg = "true";
defparam \mem~186 .power_up = "low";

dffeas \mem~218 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~218_q ),
	.prn(vcc));
defparam \mem~218 .is_wysiwyg = "true";
defparam \mem~218 .power_up = "low";

dffeas \mem~154 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~154_q ),
	.prn(vcc));
defparam \mem~154 .is_wysiwyg = "true";
defparam \mem~154 .power_up = "low";

cycloneive_lcell_comb \mem~301 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~218_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~154_q ),
	.cin(gnd),
	.combout(\mem~301_combout ),
	.cout());
defparam \mem~301 .lut_mask = 16'hFFDE;
defparam \mem~301 .sum_lutc_input = "datac";

dffeas \mem~250 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~250_q ),
	.prn(vcc));
defparam \mem~250 .is_wysiwyg = "true";
defparam \mem~250 .power_up = "low";

cycloneive_lcell_comb \mem~302 (
	.dataa(\mem~186_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~301_combout ),
	.datad(\mem~250_q ),
	.cin(gnd),
	.combout(\mem~302_combout ),
	.cout());
defparam \mem~302 .lut_mask = 16'hFFBE;
defparam \mem~302 .sum_lutc_input = "datac";

dffeas \mem~90 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~90_q ),
	.prn(vcc));
defparam \mem~90 .is_wysiwyg = "true";
defparam \mem~90 .power_up = "low";

dffeas \mem~58 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~58_q ),
	.prn(vcc));
defparam \mem~58 .is_wysiwyg = "true";
defparam \mem~58 .power_up = "low";

dffeas \mem~26 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~26_q ),
	.prn(vcc));
defparam \mem~26 .is_wysiwyg = "true";
defparam \mem~26 .power_up = "low";

cycloneive_lcell_comb \mem~303 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~58_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~26_q ),
	.cin(gnd),
	.combout(\mem~303_combout ),
	.cout());
defparam \mem~303 .lut_mask = 16'hFFDE;
defparam \mem~303 .sum_lutc_input = "datac";

dffeas \mem~122 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~122_q ),
	.prn(vcc));
defparam \mem~122 .is_wysiwyg = "true";
defparam \mem~122 .power_up = "low";

cycloneive_lcell_comb \mem~304 (
	.dataa(\mem~90_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~303_combout ),
	.datad(\mem~122_q ),
	.cin(gnd),
	.combout(\mem~304_combout ),
	.cout());
defparam \mem~304 .lut_mask = 16'hFFBE;
defparam \mem~304 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~305 (
	.dataa(\mem~302_combout ),
	.datab(\mem~304_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~305_combout ),
	.cout());
defparam \mem~305 .lut_mask = 16'hAACC;
defparam \mem~305 .sum_lutc_input = "datac";

dffeas \internal_out_payload[26] (
	.clk(clk),
	.d(\mem~305_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[26]~q ),
	.prn(vcc));
defparam \internal_out_payload[26] .is_wysiwyg = "true";
defparam \internal_out_payload[26] .power_up = "low";

dffeas \mem~171 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~171_q ),
	.prn(vcc));
defparam \mem~171 .is_wysiwyg = "true";
defparam \mem~171 .power_up = "low";

dffeas \mem~203 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~203_q ),
	.prn(vcc));
defparam \mem~203 .is_wysiwyg = "true";
defparam \mem~203 .power_up = "low";

dffeas \mem~139 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~139_q ),
	.prn(vcc));
defparam \mem~139 .is_wysiwyg = "true";
defparam \mem~139 .power_up = "low";

cycloneive_lcell_comb \mem~306 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~203_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~139_q ),
	.cin(gnd),
	.combout(\mem~306_combout ),
	.cout());
defparam \mem~306 .lut_mask = 16'hFFDE;
defparam \mem~306 .sum_lutc_input = "datac";

dffeas \mem~235 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~235_q ),
	.prn(vcc));
defparam \mem~235 .is_wysiwyg = "true";
defparam \mem~235 .power_up = "low";

cycloneive_lcell_comb \mem~307 (
	.dataa(\mem~171_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~306_combout ),
	.datad(\mem~235_q ),
	.cin(gnd),
	.combout(\mem~307_combout ),
	.cout());
defparam \mem~307 .lut_mask = 16'hFFBE;
defparam \mem~307 .sum_lutc_input = "datac";

dffeas \mem~75 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~75_q ),
	.prn(vcc));
defparam \mem~75 .is_wysiwyg = "true";
defparam \mem~75 .power_up = "low";

dffeas \mem~43 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~43_q ),
	.prn(vcc));
defparam \mem~43 .is_wysiwyg = "true";
defparam \mem~43 .power_up = "low";

dffeas \mem~11 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~11_q ),
	.prn(vcc));
defparam \mem~11 .is_wysiwyg = "true";
defparam \mem~11 .power_up = "low";

cycloneive_lcell_comb \mem~308 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~43_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~11_q ),
	.cin(gnd),
	.combout(\mem~308_combout ),
	.cout());
defparam \mem~308 .lut_mask = 16'hFFDE;
defparam \mem~308 .sum_lutc_input = "datac";

dffeas \mem~107 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~107_q ),
	.prn(vcc));
defparam \mem~107 .is_wysiwyg = "true";
defparam \mem~107 .power_up = "low";

cycloneive_lcell_comb \mem~309 (
	.dataa(\mem~75_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~308_combout ),
	.datad(\mem~107_q ),
	.cin(gnd),
	.combout(\mem~309_combout ),
	.cout());
defparam \mem~309 .lut_mask = 16'hFFBE;
defparam \mem~309 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~310 (
	.dataa(\mem~307_combout ),
	.datab(\mem~309_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~310_combout ),
	.cout());
defparam \mem~310 .lut_mask = 16'hAACC;
defparam \mem~310 .sum_lutc_input = "datac";

dffeas \internal_out_payload[11] (
	.clk(clk),
	.d(\mem~310_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[11]~q ),
	.prn(vcc));
defparam \internal_out_payload[11] .is_wysiwyg = "true";
defparam \internal_out_payload[11] .power_up = "low";

dffeas \mem~173 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~173_q ),
	.prn(vcc));
defparam \mem~173 .is_wysiwyg = "true";
defparam \mem~173 .power_up = "low";

dffeas \mem~205 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~205_q ),
	.prn(vcc));
defparam \mem~205 .is_wysiwyg = "true";
defparam \mem~205 .power_up = "low";

dffeas \mem~141 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~141_q ),
	.prn(vcc));
defparam \mem~141 .is_wysiwyg = "true";
defparam \mem~141 .power_up = "low";

cycloneive_lcell_comb \mem~311 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~205_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~141_q ),
	.cin(gnd),
	.combout(\mem~311_combout ),
	.cout());
defparam \mem~311 .lut_mask = 16'hFFDE;
defparam \mem~311 .sum_lutc_input = "datac";

dffeas \mem~237 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~237_q ),
	.prn(vcc));
defparam \mem~237 .is_wysiwyg = "true";
defparam \mem~237 .power_up = "low";

cycloneive_lcell_comb \mem~312 (
	.dataa(\mem~173_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~311_combout ),
	.datad(\mem~237_q ),
	.cin(gnd),
	.combout(\mem~312_combout ),
	.cout());
defparam \mem~312 .lut_mask = 16'hFFBE;
defparam \mem~312 .sum_lutc_input = "datac";

dffeas \mem~77 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~77_q ),
	.prn(vcc));
defparam \mem~77 .is_wysiwyg = "true";
defparam \mem~77 .power_up = "low";

dffeas \mem~45 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~45_q ),
	.prn(vcc));
defparam \mem~45 .is_wysiwyg = "true";
defparam \mem~45 .power_up = "low";

dffeas \mem~13 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~13_q ),
	.prn(vcc));
defparam \mem~13 .is_wysiwyg = "true";
defparam \mem~13 .power_up = "low";

cycloneive_lcell_comb \mem~313 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~45_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~13_q ),
	.cin(gnd),
	.combout(\mem~313_combout ),
	.cout());
defparam \mem~313 .lut_mask = 16'hFFDE;
defparam \mem~313 .sum_lutc_input = "datac";

dffeas \mem~109 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~109_q ),
	.prn(vcc));
defparam \mem~109 .is_wysiwyg = "true";
defparam \mem~109 .power_up = "low";

cycloneive_lcell_comb \mem~314 (
	.dataa(\mem~77_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~313_combout ),
	.datad(\mem~109_q ),
	.cin(gnd),
	.combout(\mem~314_combout ),
	.cout());
defparam \mem~314 .lut_mask = 16'hFFBE;
defparam \mem~314 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~315 (
	.dataa(\mem~312_combout ),
	.datab(\mem~314_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~315_combout ),
	.cout());
defparam \mem~315 .lut_mask = 16'hAACC;
defparam \mem~315 .sum_lutc_input = "datac";

dffeas \internal_out_payload[13] (
	.clk(clk),
	.d(\mem~315_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[13]~q ),
	.prn(vcc));
defparam \internal_out_payload[13] .is_wysiwyg = "true";
defparam \internal_out_payload[13] .power_up = "low";

dffeas \mem~176 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~176_q ),
	.prn(vcc));
defparam \mem~176 .is_wysiwyg = "true";
defparam \mem~176 .power_up = "low";

dffeas \mem~208 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~208_q ),
	.prn(vcc));
defparam \mem~208 .is_wysiwyg = "true";
defparam \mem~208 .power_up = "low";

dffeas \mem~144 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~144_q ),
	.prn(vcc));
defparam \mem~144 .is_wysiwyg = "true";
defparam \mem~144 .power_up = "low";

cycloneive_lcell_comb \mem~316 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~208_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~144_q ),
	.cin(gnd),
	.combout(\mem~316_combout ),
	.cout());
defparam \mem~316 .lut_mask = 16'hFFDE;
defparam \mem~316 .sum_lutc_input = "datac";

dffeas \mem~240 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~240_q ),
	.prn(vcc));
defparam \mem~240 .is_wysiwyg = "true";
defparam \mem~240 .power_up = "low";

cycloneive_lcell_comb \mem~317 (
	.dataa(\mem~176_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~316_combout ),
	.datad(\mem~240_q ),
	.cin(gnd),
	.combout(\mem~317_combout ),
	.cout());
defparam \mem~317 .lut_mask = 16'hFFBE;
defparam \mem~317 .sum_lutc_input = "datac";

dffeas \mem~80 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~80_q ),
	.prn(vcc));
defparam \mem~80 .is_wysiwyg = "true";
defparam \mem~80 .power_up = "low";

dffeas \mem~48 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~48_q ),
	.prn(vcc));
defparam \mem~48 .is_wysiwyg = "true";
defparam \mem~48 .power_up = "low";

dffeas \mem~16 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~16_q ),
	.prn(vcc));
defparam \mem~16 .is_wysiwyg = "true";
defparam \mem~16 .power_up = "low";

cycloneive_lcell_comb \mem~318 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~48_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~16_q ),
	.cin(gnd),
	.combout(\mem~318_combout ),
	.cout());
defparam \mem~318 .lut_mask = 16'hFFDE;
defparam \mem~318 .sum_lutc_input = "datac";

dffeas \mem~112 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~112_q ),
	.prn(vcc));
defparam \mem~112 .is_wysiwyg = "true";
defparam \mem~112 .power_up = "low";

cycloneive_lcell_comb \mem~319 (
	.dataa(\mem~80_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~318_combout ),
	.datad(\mem~112_q ),
	.cin(gnd),
	.combout(\mem~319_combout ),
	.cout());
defparam \mem~319 .lut_mask = 16'hFFBE;
defparam \mem~319 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~320 (
	.dataa(\mem~317_combout ),
	.datab(\mem~319_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~320_combout ),
	.cout());
defparam \mem~320 .lut_mask = 16'hAACC;
defparam \mem~320 .sum_lutc_input = "datac";

dffeas \internal_out_payload[16] (
	.clk(clk),
	.d(\mem~320_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[16]~q ),
	.prn(vcc));
defparam \internal_out_payload[16] .is_wysiwyg = "true";
defparam \internal_out_payload[16] .power_up = "low";

dffeas \mem~172 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~172_q ),
	.prn(vcc));
defparam \mem~172 .is_wysiwyg = "true";
defparam \mem~172 .power_up = "low";

dffeas \mem~204 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~204_q ),
	.prn(vcc));
defparam \mem~204 .is_wysiwyg = "true";
defparam \mem~204 .power_up = "low";

dffeas \mem~140 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~140_q ),
	.prn(vcc));
defparam \mem~140 .is_wysiwyg = "true";
defparam \mem~140 .power_up = "low";

cycloneive_lcell_comb \mem~321 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~204_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~140_q ),
	.cin(gnd),
	.combout(\mem~321_combout ),
	.cout());
defparam \mem~321 .lut_mask = 16'hFFDE;
defparam \mem~321 .sum_lutc_input = "datac";

dffeas \mem~236 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~236_q ),
	.prn(vcc));
defparam \mem~236 .is_wysiwyg = "true";
defparam \mem~236 .power_up = "low";

cycloneive_lcell_comb \mem~322 (
	.dataa(\mem~172_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~321_combout ),
	.datad(\mem~236_q ),
	.cin(gnd),
	.combout(\mem~322_combout ),
	.cout());
defparam \mem~322 .lut_mask = 16'hFFBE;
defparam \mem~322 .sum_lutc_input = "datac";

dffeas \mem~76 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~76_q ),
	.prn(vcc));
defparam \mem~76 .is_wysiwyg = "true";
defparam \mem~76 .power_up = "low";

dffeas \mem~44 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~44_q ),
	.prn(vcc));
defparam \mem~44 .is_wysiwyg = "true";
defparam \mem~44 .power_up = "low";

dffeas \mem~12 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~12_q ),
	.prn(vcc));
defparam \mem~12 .is_wysiwyg = "true";
defparam \mem~12 .power_up = "low";

cycloneive_lcell_comb \mem~323 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~44_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~12_q ),
	.cin(gnd),
	.combout(\mem~323_combout ),
	.cout());
defparam \mem~323 .lut_mask = 16'hFFDE;
defparam \mem~323 .sum_lutc_input = "datac";

dffeas \mem~108 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~108_q ),
	.prn(vcc));
defparam \mem~108 .is_wysiwyg = "true";
defparam \mem~108 .power_up = "low";

cycloneive_lcell_comb \mem~324 (
	.dataa(\mem~76_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~323_combout ),
	.datad(\mem~108_q ),
	.cin(gnd),
	.combout(\mem~324_combout ),
	.cout());
defparam \mem~324 .lut_mask = 16'hFFBE;
defparam \mem~324 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~325 (
	.dataa(\mem~322_combout ),
	.datab(\mem~324_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~325_combout ),
	.cout());
defparam \mem~325 .lut_mask = 16'hAACC;
defparam \mem~325 .sum_lutc_input = "datac";

dffeas \internal_out_payload[12] (
	.clk(clk),
	.d(\mem~325_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[12]~q ),
	.prn(vcc));
defparam \internal_out_payload[12] .is_wysiwyg = "true";
defparam \internal_out_payload[12] .power_up = "low";

dffeas \mem~165 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~165_q ),
	.prn(vcc));
defparam \mem~165 .is_wysiwyg = "true";
defparam \mem~165 .power_up = "low";

dffeas \mem~197 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~197_q ),
	.prn(vcc));
defparam \mem~197 .is_wysiwyg = "true";
defparam \mem~197 .power_up = "low";

dffeas \mem~133 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~133_q ),
	.prn(vcc));
defparam \mem~133 .is_wysiwyg = "true";
defparam \mem~133 .power_up = "low";

cycloneive_lcell_comb \mem~326 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~197_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~133_q ),
	.cin(gnd),
	.combout(\mem~326_combout ),
	.cout());
defparam \mem~326 .lut_mask = 16'hFFDE;
defparam \mem~326 .sum_lutc_input = "datac";

dffeas \mem~229 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~229_q ),
	.prn(vcc));
defparam \mem~229 .is_wysiwyg = "true";
defparam \mem~229 .power_up = "low";

cycloneive_lcell_comb \mem~327 (
	.dataa(\mem~165_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~326_combout ),
	.datad(\mem~229_q ),
	.cin(gnd),
	.combout(\mem~327_combout ),
	.cout());
defparam \mem~327 .lut_mask = 16'hFFBE;
defparam \mem~327 .sum_lutc_input = "datac";

dffeas \mem~69 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~69_q ),
	.prn(vcc));
defparam \mem~69 .is_wysiwyg = "true";
defparam \mem~69 .power_up = "low";

dffeas \mem~37 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~37_q ),
	.prn(vcc));
defparam \mem~37 .is_wysiwyg = "true";
defparam \mem~37 .power_up = "low";

dffeas \mem~5 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~5_q ),
	.prn(vcc));
defparam \mem~5 .is_wysiwyg = "true";
defparam \mem~5 .power_up = "low";

cycloneive_lcell_comb \mem~328 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~37_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~5_q ),
	.cin(gnd),
	.combout(\mem~328_combout ),
	.cout());
defparam \mem~328 .lut_mask = 16'hFFDE;
defparam \mem~328 .sum_lutc_input = "datac";

dffeas \mem~101 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~101_q ),
	.prn(vcc));
defparam \mem~101 .is_wysiwyg = "true";
defparam \mem~101 .power_up = "low";

cycloneive_lcell_comb \mem~329 (
	.dataa(\mem~69_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~328_combout ),
	.datad(\mem~101_q ),
	.cin(gnd),
	.combout(\mem~329_combout ),
	.cout());
defparam \mem~329 .lut_mask = 16'hFFBE;
defparam \mem~329 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~330 (
	.dataa(\mem~327_combout ),
	.datab(\mem~329_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~330_combout ),
	.cout());
defparam \mem~330 .lut_mask = 16'hAACC;
defparam \mem~330 .sum_lutc_input = "datac";

dffeas \internal_out_payload[5] (
	.clk(clk),
	.d(\mem~330_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[5]~q ),
	.prn(vcc));
defparam \internal_out_payload[5] .is_wysiwyg = "true";
defparam \internal_out_payload[5] .power_up = "low";

dffeas \mem~174 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~174_q ),
	.prn(vcc));
defparam \mem~174 .is_wysiwyg = "true";
defparam \mem~174 .power_up = "low";

dffeas \mem~206 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~206_q ),
	.prn(vcc));
defparam \mem~206 .is_wysiwyg = "true";
defparam \mem~206 .power_up = "low";

dffeas \mem~142 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~142_q ),
	.prn(vcc));
defparam \mem~142 .is_wysiwyg = "true";
defparam \mem~142 .power_up = "low";

cycloneive_lcell_comb \mem~331 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~206_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~142_q ),
	.cin(gnd),
	.combout(\mem~331_combout ),
	.cout());
defparam \mem~331 .lut_mask = 16'hFFDE;
defparam \mem~331 .sum_lutc_input = "datac";

dffeas \mem~238 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~238_q ),
	.prn(vcc));
defparam \mem~238 .is_wysiwyg = "true";
defparam \mem~238 .power_up = "low";

cycloneive_lcell_comb \mem~332 (
	.dataa(\mem~174_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~331_combout ),
	.datad(\mem~238_q ),
	.cin(gnd),
	.combout(\mem~332_combout ),
	.cout());
defparam \mem~332 .lut_mask = 16'hFFBE;
defparam \mem~332 .sum_lutc_input = "datac";

dffeas \mem~78 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~78_q ),
	.prn(vcc));
defparam \mem~78 .is_wysiwyg = "true";
defparam \mem~78 .power_up = "low";

dffeas \mem~46 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~46_q ),
	.prn(vcc));
defparam \mem~46 .is_wysiwyg = "true";
defparam \mem~46 .power_up = "low";

dffeas \mem~14 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~14_q ),
	.prn(vcc));
defparam \mem~14 .is_wysiwyg = "true";
defparam \mem~14 .power_up = "low";

cycloneive_lcell_comb \mem~333 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~46_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~14_q ),
	.cin(gnd),
	.combout(\mem~333_combout ),
	.cout());
defparam \mem~333 .lut_mask = 16'hFFDE;
defparam \mem~333 .sum_lutc_input = "datac";

dffeas \mem~110 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~110_q ),
	.prn(vcc));
defparam \mem~110 .is_wysiwyg = "true";
defparam \mem~110 .power_up = "low";

cycloneive_lcell_comb \mem~334 (
	.dataa(\mem~78_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~333_combout ),
	.datad(\mem~110_q ),
	.cin(gnd),
	.combout(\mem~334_combout ),
	.cout());
defparam \mem~334 .lut_mask = 16'hFFBE;
defparam \mem~334 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~335 (
	.dataa(\mem~332_combout ),
	.datab(\mem~334_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~335_combout ),
	.cout());
defparam \mem~335 .lut_mask = 16'hAACC;
defparam \mem~335 .sum_lutc_input = "datac";

dffeas \internal_out_payload[14] (
	.clk(clk),
	.d(\mem~335_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[14]~q ),
	.prn(vcc));
defparam \internal_out_payload[14] .is_wysiwyg = "true";
defparam \internal_out_payload[14] .power_up = "low";

dffeas \mem~175 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~175_q ),
	.prn(vcc));
defparam \mem~175 .is_wysiwyg = "true";
defparam \mem~175 .power_up = "low";

dffeas \mem~207 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~207_q ),
	.prn(vcc));
defparam \mem~207 .is_wysiwyg = "true";
defparam \mem~207 .power_up = "low";

dffeas \mem~143 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~143_q ),
	.prn(vcc));
defparam \mem~143 .is_wysiwyg = "true";
defparam \mem~143 .power_up = "low";

cycloneive_lcell_comb \mem~336 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~207_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~143_q ),
	.cin(gnd),
	.combout(\mem~336_combout ),
	.cout());
defparam \mem~336 .lut_mask = 16'hFFDE;
defparam \mem~336 .sum_lutc_input = "datac";

dffeas \mem~239 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~239_q ),
	.prn(vcc));
defparam \mem~239 .is_wysiwyg = "true";
defparam \mem~239 .power_up = "low";

cycloneive_lcell_comb \mem~337 (
	.dataa(\mem~175_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~336_combout ),
	.datad(\mem~239_q ),
	.cin(gnd),
	.combout(\mem~337_combout ),
	.cout());
defparam \mem~337 .lut_mask = 16'hFFBE;
defparam \mem~337 .sum_lutc_input = "datac";

dffeas \mem~79 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~79_q ),
	.prn(vcc));
defparam \mem~79 .is_wysiwyg = "true";
defparam \mem~79 .power_up = "low";

dffeas \mem~47 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~47_q ),
	.prn(vcc));
defparam \mem~47 .is_wysiwyg = "true";
defparam \mem~47 .power_up = "low";

dffeas \mem~15 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~15_q ),
	.prn(vcc));
defparam \mem~15 .is_wysiwyg = "true";
defparam \mem~15 .power_up = "low";

cycloneive_lcell_comb \mem~338 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~47_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~15_q ),
	.cin(gnd),
	.combout(\mem~338_combout ),
	.cout());
defparam \mem~338 .lut_mask = 16'hFFDE;
defparam \mem~338 .sum_lutc_input = "datac";

dffeas \mem~111 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~111_q ),
	.prn(vcc));
defparam \mem~111 .is_wysiwyg = "true";
defparam \mem~111 .power_up = "low";

cycloneive_lcell_comb \mem~339 (
	.dataa(\mem~79_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~338_combout ),
	.datad(\mem~111_q ),
	.cin(gnd),
	.combout(\mem~339_combout ),
	.cout());
defparam \mem~339 .lut_mask = 16'hFFBE;
defparam \mem~339 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~340 (
	.dataa(\mem~337_combout ),
	.datab(\mem~339_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~340_combout ),
	.cout());
defparam \mem~340 .lut_mask = 16'hAACC;
defparam \mem~340 .sum_lutc_input = "datac";

dffeas \internal_out_payload[15] (
	.clk(clk),
	.d(\mem~340_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[15]~q ),
	.prn(vcc));
defparam \internal_out_payload[15] .is_wysiwyg = "true";
defparam \internal_out_payload[15] .power_up = "low";

dffeas \mem~170 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~170_q ),
	.prn(vcc));
defparam \mem~170 .is_wysiwyg = "true";
defparam \mem~170 .power_up = "low";

dffeas \mem~202 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~202_q ),
	.prn(vcc));
defparam \mem~202 .is_wysiwyg = "true";
defparam \mem~202 .power_up = "low";

dffeas \mem~138 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~138_q ),
	.prn(vcc));
defparam \mem~138 .is_wysiwyg = "true";
defparam \mem~138 .power_up = "low";

cycloneive_lcell_comb \mem~341 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~202_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~138_q ),
	.cin(gnd),
	.combout(\mem~341_combout ),
	.cout());
defparam \mem~341 .lut_mask = 16'hFFDE;
defparam \mem~341 .sum_lutc_input = "datac";

dffeas \mem~234 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~234_q ),
	.prn(vcc));
defparam \mem~234 .is_wysiwyg = "true";
defparam \mem~234 .power_up = "low";

cycloneive_lcell_comb \mem~342 (
	.dataa(\mem~170_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~341_combout ),
	.datad(\mem~234_q ),
	.cin(gnd),
	.combout(\mem~342_combout ),
	.cout());
defparam \mem~342 .lut_mask = 16'hFFBE;
defparam \mem~342 .sum_lutc_input = "datac";

dffeas \mem~74 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~74_q ),
	.prn(vcc));
defparam \mem~74 .is_wysiwyg = "true";
defparam \mem~74 .power_up = "low";

dffeas \mem~42 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~42_q ),
	.prn(vcc));
defparam \mem~42 .is_wysiwyg = "true";
defparam \mem~42 .power_up = "low";

dffeas \mem~10 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~10_q ),
	.prn(vcc));
defparam \mem~10 .is_wysiwyg = "true";
defparam \mem~10 .power_up = "low";

cycloneive_lcell_comb \mem~343 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~42_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~10_q ),
	.cin(gnd),
	.combout(\mem~343_combout ),
	.cout());
defparam \mem~343 .lut_mask = 16'hFFDE;
defparam \mem~343 .sum_lutc_input = "datac";

dffeas \mem~106 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~106_q ),
	.prn(vcc));
defparam \mem~106 .is_wysiwyg = "true";
defparam \mem~106 .power_up = "low";

cycloneive_lcell_comb \mem~344 (
	.dataa(\mem~74_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~343_combout ),
	.datad(\mem~106_q ),
	.cin(gnd),
	.combout(\mem~344_combout ),
	.cout());
defparam \mem~344 .lut_mask = 16'hFFBE;
defparam \mem~344 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~345 (
	.dataa(\mem~342_combout ),
	.datab(\mem~344_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~345_combout ),
	.cout());
defparam \mem~345 .lut_mask = 16'hAACC;
defparam \mem~345 .sum_lutc_input = "datac";

dffeas \internal_out_payload[10] (
	.clk(clk),
	.d(\mem~345_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[10]~q ),
	.prn(vcc));
defparam \internal_out_payload[10] .is_wysiwyg = "true";
defparam \internal_out_payload[10] .power_up = "low";

dffeas \mem~169 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~169_q ),
	.prn(vcc));
defparam \mem~169 .is_wysiwyg = "true";
defparam \mem~169 .power_up = "low";

dffeas \mem~201 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~201_q ),
	.prn(vcc));
defparam \mem~201 .is_wysiwyg = "true";
defparam \mem~201 .power_up = "low";

dffeas \mem~137 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~137_q ),
	.prn(vcc));
defparam \mem~137 .is_wysiwyg = "true";
defparam \mem~137 .power_up = "low";

cycloneive_lcell_comb \mem~346 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~201_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~137_q ),
	.cin(gnd),
	.combout(\mem~346_combout ),
	.cout());
defparam \mem~346 .lut_mask = 16'hFFDE;
defparam \mem~346 .sum_lutc_input = "datac";

dffeas \mem~233 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~233_q ),
	.prn(vcc));
defparam \mem~233 .is_wysiwyg = "true";
defparam \mem~233 .power_up = "low";

cycloneive_lcell_comb \mem~347 (
	.dataa(\mem~169_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~346_combout ),
	.datad(\mem~233_q ),
	.cin(gnd),
	.combout(\mem~347_combout ),
	.cout());
defparam \mem~347 .lut_mask = 16'hFFBE;
defparam \mem~347 .sum_lutc_input = "datac";

dffeas \mem~73 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~73_q ),
	.prn(vcc));
defparam \mem~73 .is_wysiwyg = "true";
defparam \mem~73 .power_up = "low";

dffeas \mem~41 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~41_q ),
	.prn(vcc));
defparam \mem~41 .is_wysiwyg = "true";
defparam \mem~41 .power_up = "low";

dffeas \mem~9 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~9_q ),
	.prn(vcc));
defparam \mem~9 .is_wysiwyg = "true";
defparam \mem~9 .power_up = "low";

cycloneive_lcell_comb \mem~348 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~41_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~9_q ),
	.cin(gnd),
	.combout(\mem~348_combout ),
	.cout());
defparam \mem~348 .lut_mask = 16'hFFDE;
defparam \mem~348 .sum_lutc_input = "datac";

dffeas \mem~105 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~105_q ),
	.prn(vcc));
defparam \mem~105 .is_wysiwyg = "true";
defparam \mem~105 .power_up = "low";

cycloneive_lcell_comb \mem~349 (
	.dataa(\mem~73_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~348_combout ),
	.datad(\mem~105_q ),
	.cin(gnd),
	.combout(\mem~349_combout ),
	.cout());
defparam \mem~349 .lut_mask = 16'hFFBE;
defparam \mem~349 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~350 (
	.dataa(\mem~347_combout ),
	.datab(\mem~349_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~350_combout ),
	.cout());
defparam \mem~350 .lut_mask = 16'hAACC;
defparam \mem~350 .sum_lutc_input = "datac";

dffeas \internal_out_payload[9] (
	.clk(clk),
	.d(\mem~350_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[9]~q ),
	.prn(vcc));
defparam \internal_out_payload[9] .is_wysiwyg = "true";
defparam \internal_out_payload[9] .power_up = "low";

dffeas \mem~168 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~168_q ),
	.prn(vcc));
defparam \mem~168 .is_wysiwyg = "true";
defparam \mem~168 .power_up = "low";

dffeas \mem~200 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~200_q ),
	.prn(vcc));
defparam \mem~200 .is_wysiwyg = "true";
defparam \mem~200 .power_up = "low";

dffeas \mem~136 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~136_q ),
	.prn(vcc));
defparam \mem~136 .is_wysiwyg = "true";
defparam \mem~136 .power_up = "low";

cycloneive_lcell_comb \mem~351 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~200_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~136_q ),
	.cin(gnd),
	.combout(\mem~351_combout ),
	.cout());
defparam \mem~351 .lut_mask = 16'hFFDE;
defparam \mem~351 .sum_lutc_input = "datac";

dffeas \mem~232 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~232_q ),
	.prn(vcc));
defparam \mem~232 .is_wysiwyg = "true";
defparam \mem~232 .power_up = "low";

cycloneive_lcell_comb \mem~352 (
	.dataa(\mem~168_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~351_combout ),
	.datad(\mem~232_q ),
	.cin(gnd),
	.combout(\mem~352_combout ),
	.cout());
defparam \mem~352 .lut_mask = 16'hFFBE;
defparam \mem~352 .sum_lutc_input = "datac";

dffeas \mem~72 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~72_q ),
	.prn(vcc));
defparam \mem~72 .is_wysiwyg = "true";
defparam \mem~72 .power_up = "low";

dffeas \mem~40 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~40_q ),
	.prn(vcc));
defparam \mem~40 .is_wysiwyg = "true";
defparam \mem~40 .power_up = "low";

dffeas \mem~8 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~8_q ),
	.prn(vcc));
defparam \mem~8 .is_wysiwyg = "true";
defparam \mem~8 .power_up = "low";

cycloneive_lcell_comb \mem~353 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~40_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~8_q ),
	.cin(gnd),
	.combout(\mem~353_combout ),
	.cout());
defparam \mem~353 .lut_mask = 16'hFFDE;
defparam \mem~353 .sum_lutc_input = "datac";

dffeas \mem~104 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~104_q ),
	.prn(vcc));
defparam \mem~104 .is_wysiwyg = "true";
defparam \mem~104 .power_up = "low";

cycloneive_lcell_comb \mem~354 (
	.dataa(\mem~72_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~353_combout ),
	.datad(\mem~104_q ),
	.cin(gnd),
	.combout(\mem~354_combout ),
	.cout());
defparam \mem~354 .lut_mask = 16'hFFBE;
defparam \mem~354 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~355 (
	.dataa(\mem~352_combout ),
	.datab(\mem~354_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~355_combout ),
	.cout());
defparam \mem~355 .lut_mask = 16'hAACC;
defparam \mem~355 .sum_lutc_input = "datac";

dffeas \internal_out_payload[8] (
	.clk(clk),
	.d(\mem~355_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[8]~q ),
	.prn(vcc));
defparam \internal_out_payload[8] .is_wysiwyg = "true";
defparam \internal_out_payload[8] .power_up = "low";

dffeas \mem~167 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~167_q ),
	.prn(vcc));
defparam \mem~167 .is_wysiwyg = "true";
defparam \mem~167 .power_up = "low";

dffeas \mem~199 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~199_q ),
	.prn(vcc));
defparam \mem~199 .is_wysiwyg = "true";
defparam \mem~199 .power_up = "low";

dffeas \mem~135 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~135_q ),
	.prn(vcc));
defparam \mem~135 .is_wysiwyg = "true";
defparam \mem~135 .power_up = "low";

cycloneive_lcell_comb \mem~356 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~199_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~135_q ),
	.cin(gnd),
	.combout(\mem~356_combout ),
	.cout());
defparam \mem~356 .lut_mask = 16'hFFDE;
defparam \mem~356 .sum_lutc_input = "datac";

dffeas \mem~231 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~231_q ),
	.prn(vcc));
defparam \mem~231 .is_wysiwyg = "true";
defparam \mem~231 .power_up = "low";

cycloneive_lcell_comb \mem~357 (
	.dataa(\mem~167_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~356_combout ),
	.datad(\mem~231_q ),
	.cin(gnd),
	.combout(\mem~357_combout ),
	.cout());
defparam \mem~357 .lut_mask = 16'hFFBE;
defparam \mem~357 .sum_lutc_input = "datac";

dffeas \mem~71 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~71_q ),
	.prn(vcc));
defparam \mem~71 .is_wysiwyg = "true";
defparam \mem~71 .power_up = "low";

dffeas \mem~39 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~39_q ),
	.prn(vcc));
defparam \mem~39 .is_wysiwyg = "true";
defparam \mem~39 .power_up = "low";

dffeas \mem~7 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~7_q ),
	.prn(vcc));
defparam \mem~7 .is_wysiwyg = "true";
defparam \mem~7 .power_up = "low";

cycloneive_lcell_comb \mem~358 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~39_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~7_q ),
	.cin(gnd),
	.combout(\mem~358_combout ),
	.cout());
defparam \mem~358 .lut_mask = 16'hFFDE;
defparam \mem~358 .sum_lutc_input = "datac";

dffeas \mem~103 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~103_q ),
	.prn(vcc));
defparam \mem~103 .is_wysiwyg = "true";
defparam \mem~103 .power_up = "low";

cycloneive_lcell_comb \mem~359 (
	.dataa(\mem~71_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~358_combout ),
	.datad(\mem~103_q ),
	.cin(gnd),
	.combout(\mem~359_combout ),
	.cout());
defparam \mem~359 .lut_mask = 16'hFFBE;
defparam \mem~359 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~360 (
	.dataa(\mem~357_combout ),
	.datab(\mem~359_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~360_combout ),
	.cout());
defparam \mem~360 .lut_mask = 16'hAACC;
defparam \mem~360 .sum_lutc_input = "datac";

dffeas \internal_out_payload[7] (
	.clk(clk),
	.d(\mem~360_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[7]~q ),
	.prn(vcc));
defparam \internal_out_payload[7] .is_wysiwyg = "true";
defparam \internal_out_payload[7] .power_up = "low";

dffeas \mem~166 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~166_q ),
	.prn(vcc));
defparam \mem~166 .is_wysiwyg = "true";
defparam \mem~166 .power_up = "low";

dffeas \mem~198 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~198_q ),
	.prn(vcc));
defparam \mem~198 .is_wysiwyg = "true";
defparam \mem~198 .power_up = "low";

dffeas \mem~134 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~134_q ),
	.prn(vcc));
defparam \mem~134 .is_wysiwyg = "true";
defparam \mem~134 .power_up = "low";

cycloneive_lcell_comb \mem~361 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~198_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~134_q ),
	.cin(gnd),
	.combout(\mem~361_combout ),
	.cout());
defparam \mem~361 .lut_mask = 16'hFFDE;
defparam \mem~361 .sum_lutc_input = "datac";

dffeas \mem~230 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~230_q ),
	.prn(vcc));
defparam \mem~230 .is_wysiwyg = "true";
defparam \mem~230 .power_up = "low";

cycloneive_lcell_comb \mem~362 (
	.dataa(\mem~166_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~361_combout ),
	.datad(\mem~230_q ),
	.cin(gnd),
	.combout(\mem~362_combout ),
	.cout());
defparam \mem~362 .lut_mask = 16'hFFBE;
defparam \mem~362 .sum_lutc_input = "datac";

dffeas \mem~70 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~70_q ),
	.prn(vcc));
defparam \mem~70 .is_wysiwyg = "true";
defparam \mem~70 .power_up = "low";

dffeas \mem~38 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~38_q ),
	.prn(vcc));
defparam \mem~38 .is_wysiwyg = "true";
defparam \mem~38 .power_up = "low";

dffeas \mem~6 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~6_q ),
	.prn(vcc));
defparam \mem~6 .is_wysiwyg = "true";
defparam \mem~6 .power_up = "low";

cycloneive_lcell_comb \mem~363 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~38_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~6_q ),
	.cin(gnd),
	.combout(\mem~363_combout ),
	.cout());
defparam \mem~363 .lut_mask = 16'hFFDE;
defparam \mem~363 .sum_lutc_input = "datac";

dffeas \mem~102 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~102_q ),
	.prn(vcc));
defparam \mem~102 .is_wysiwyg = "true";
defparam \mem~102 .power_up = "low";

cycloneive_lcell_comb \mem~364 (
	.dataa(\mem~70_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~363_combout ),
	.datad(\mem~102_q ),
	.cin(gnd),
	.combout(\mem~364_combout ),
	.cout());
defparam \mem~364 .lut_mask = 16'hFFBE;
defparam \mem~364 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~365 (
	.dataa(\mem~362_combout ),
	.datab(\mem~364_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~365_combout ),
	.cout());
defparam \mem~365 .lut_mask = 16'hAACC;
defparam \mem~365 .sum_lutc_input = "datac";

dffeas \internal_out_payload[6] (
	.clk(clk),
	.d(\mem~365_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[6]~q ),
	.prn(vcc));
defparam \internal_out_payload[6] .is_wysiwyg = "true";
defparam \internal_out_payload[6] .power_up = "low";

dffeas \mem~180 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~180_q ),
	.prn(vcc));
defparam \mem~180 .is_wysiwyg = "true";
defparam \mem~180 .power_up = "low";

dffeas \mem~212 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~212_q ),
	.prn(vcc));
defparam \mem~212 .is_wysiwyg = "true";
defparam \mem~212 .power_up = "low";

dffeas \mem~148 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~148_q ),
	.prn(vcc));
defparam \mem~148 .is_wysiwyg = "true";
defparam \mem~148 .power_up = "low";

cycloneive_lcell_comb \mem~366 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~212_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~148_q ),
	.cin(gnd),
	.combout(\mem~366_combout ),
	.cout());
defparam \mem~366 .lut_mask = 16'hFFDE;
defparam \mem~366 .sum_lutc_input = "datac";

dffeas \mem~244 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~244_q ),
	.prn(vcc));
defparam \mem~244 .is_wysiwyg = "true";
defparam \mem~244 .power_up = "low";

cycloneive_lcell_comb \mem~367 (
	.dataa(\mem~180_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~366_combout ),
	.datad(\mem~244_q ),
	.cin(gnd),
	.combout(\mem~367_combout ),
	.cout());
defparam \mem~367 .lut_mask = 16'hFFBE;
defparam \mem~367 .sum_lutc_input = "datac";

dffeas \mem~84 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~84_q ),
	.prn(vcc));
defparam \mem~84 .is_wysiwyg = "true";
defparam \mem~84 .power_up = "low";

dffeas \mem~52 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~52_q ),
	.prn(vcc));
defparam \mem~52 .is_wysiwyg = "true";
defparam \mem~52 .power_up = "low";

dffeas \mem~20 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~20_q ),
	.prn(vcc));
defparam \mem~20 .is_wysiwyg = "true";
defparam \mem~20 .power_up = "low";

cycloneive_lcell_comb \mem~368 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~52_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~20_q ),
	.cin(gnd),
	.combout(\mem~368_combout ),
	.cout());
defparam \mem~368 .lut_mask = 16'hFFDE;
defparam \mem~368 .sum_lutc_input = "datac";

dffeas \mem~116 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~116_q ),
	.prn(vcc));
defparam \mem~116 .is_wysiwyg = "true";
defparam \mem~116 .power_up = "low";

cycloneive_lcell_comb \mem~369 (
	.dataa(\mem~84_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~368_combout ),
	.datad(\mem~116_q ),
	.cin(gnd),
	.combout(\mem~369_combout ),
	.cout());
defparam \mem~369 .lut_mask = 16'hFFBE;
defparam \mem~369 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~370 (
	.dataa(\mem~367_combout ),
	.datab(\mem~369_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~370_combout ),
	.cout());
defparam \mem~370 .lut_mask = 16'hAACC;
defparam \mem~370 .sum_lutc_input = "datac";

dffeas \internal_out_payload[20] (
	.clk(clk),
	.d(\mem~370_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[20]~q ),
	.prn(vcc));
defparam \internal_out_payload[20] .is_wysiwyg = "true";
defparam \internal_out_payload[20] .power_up = "low";

dffeas \mem~178 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~178_q ),
	.prn(vcc));
defparam \mem~178 .is_wysiwyg = "true";
defparam \mem~178 .power_up = "low";

dffeas \mem~210 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~210_q ),
	.prn(vcc));
defparam \mem~210 .is_wysiwyg = "true";
defparam \mem~210 .power_up = "low";

dffeas \mem~146 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~146_q ),
	.prn(vcc));
defparam \mem~146 .is_wysiwyg = "true";
defparam \mem~146 .power_up = "low";

cycloneive_lcell_comb \mem~371 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~210_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~146_q ),
	.cin(gnd),
	.combout(\mem~371_combout ),
	.cout());
defparam \mem~371 .lut_mask = 16'hFFDE;
defparam \mem~371 .sum_lutc_input = "datac";

dffeas \mem~242 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~242_q ),
	.prn(vcc));
defparam \mem~242 .is_wysiwyg = "true";
defparam \mem~242 .power_up = "low";

cycloneive_lcell_comb \mem~372 (
	.dataa(\mem~178_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~371_combout ),
	.datad(\mem~242_q ),
	.cin(gnd),
	.combout(\mem~372_combout ),
	.cout());
defparam \mem~372 .lut_mask = 16'hFFBE;
defparam \mem~372 .sum_lutc_input = "datac";

dffeas \mem~82 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~82_q ),
	.prn(vcc));
defparam \mem~82 .is_wysiwyg = "true";
defparam \mem~82 .power_up = "low";

dffeas \mem~50 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~50_q ),
	.prn(vcc));
defparam \mem~50 .is_wysiwyg = "true";
defparam \mem~50 .power_up = "low";

dffeas \mem~18 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~18_q ),
	.prn(vcc));
defparam \mem~18 .is_wysiwyg = "true";
defparam \mem~18 .power_up = "low";

cycloneive_lcell_comb \mem~373 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~50_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~18_q ),
	.cin(gnd),
	.combout(\mem~373_combout ),
	.cout());
defparam \mem~373 .lut_mask = 16'hFFDE;
defparam \mem~373 .sum_lutc_input = "datac";

dffeas \mem~114 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~114_q ),
	.prn(vcc));
defparam \mem~114 .is_wysiwyg = "true";
defparam \mem~114 .power_up = "low";

cycloneive_lcell_comb \mem~374 (
	.dataa(\mem~82_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~373_combout ),
	.datad(\mem~114_q ),
	.cin(gnd),
	.combout(\mem~374_combout ),
	.cout());
defparam \mem~374 .lut_mask = 16'hFFBE;
defparam \mem~374 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~375 (
	.dataa(\mem~372_combout ),
	.datab(\mem~374_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~375_combout ),
	.cout());
defparam \mem~375 .lut_mask = 16'hAACC;
defparam \mem~375 .sum_lutc_input = "datac";

dffeas \internal_out_payload[18] (
	.clk(clk),
	.d(\mem~375_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[18]~q ),
	.prn(vcc));
defparam \internal_out_payload[18] .is_wysiwyg = "true";
defparam \internal_out_payload[18] .power_up = "low";

dffeas \mem~179 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~179_q ),
	.prn(vcc));
defparam \mem~179 .is_wysiwyg = "true";
defparam \mem~179 .power_up = "low";

dffeas \mem~211 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~211_q ),
	.prn(vcc));
defparam \mem~211 .is_wysiwyg = "true";
defparam \mem~211 .power_up = "low";

dffeas \mem~147 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~147_q ),
	.prn(vcc));
defparam \mem~147 .is_wysiwyg = "true";
defparam \mem~147 .power_up = "low";

cycloneive_lcell_comb \mem~376 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~211_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~147_q ),
	.cin(gnd),
	.combout(\mem~376_combout ),
	.cout());
defparam \mem~376 .lut_mask = 16'hFFDE;
defparam \mem~376 .sum_lutc_input = "datac";

dffeas \mem~243 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~243_q ),
	.prn(vcc));
defparam \mem~243 .is_wysiwyg = "true";
defparam \mem~243 .power_up = "low";

cycloneive_lcell_comb \mem~377 (
	.dataa(\mem~179_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~376_combout ),
	.datad(\mem~243_q ),
	.cin(gnd),
	.combout(\mem~377_combout ),
	.cout());
defparam \mem~377 .lut_mask = 16'hFFBE;
defparam \mem~377 .sum_lutc_input = "datac";

dffeas \mem~83 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~83_q ),
	.prn(vcc));
defparam \mem~83 .is_wysiwyg = "true";
defparam \mem~83 .power_up = "low";

dffeas \mem~51 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~51_q ),
	.prn(vcc));
defparam \mem~51 .is_wysiwyg = "true";
defparam \mem~51 .power_up = "low";

dffeas \mem~19 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~19_q ),
	.prn(vcc));
defparam \mem~19 .is_wysiwyg = "true";
defparam \mem~19 .power_up = "low";

cycloneive_lcell_comb \mem~378 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~51_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~19_q ),
	.cin(gnd),
	.combout(\mem~378_combout ),
	.cout());
defparam \mem~378 .lut_mask = 16'hFFDE;
defparam \mem~378 .sum_lutc_input = "datac";

dffeas \mem~115 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~115_q ),
	.prn(vcc));
defparam \mem~115 .is_wysiwyg = "true";
defparam \mem~115 .power_up = "low";

cycloneive_lcell_comb \mem~379 (
	.dataa(\mem~83_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~378_combout ),
	.datad(\mem~115_q ),
	.cin(gnd),
	.combout(\mem~379_combout ),
	.cout());
defparam \mem~379 .lut_mask = 16'hFFBE;
defparam \mem~379 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~380 (
	.dataa(\mem~377_combout ),
	.datab(\mem~379_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~380_combout ),
	.cout());
defparam \mem~380 .lut_mask = 16'hAACC;
defparam \mem~380 .sum_lutc_input = "datac";

dffeas \internal_out_payload[19] (
	.clk(clk),
	.d(\mem~380_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[19]~q ),
	.prn(vcc));
defparam \internal_out_payload[19] .is_wysiwyg = "true";
defparam \internal_out_payload[19] .power_up = "low";

dffeas \mem~177 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~177_q ),
	.prn(vcc));
defparam \mem~177 .is_wysiwyg = "true";
defparam \mem~177 .power_up = "low";

dffeas \mem~209 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~209_q ),
	.prn(vcc));
defparam \mem~209 .is_wysiwyg = "true";
defparam \mem~209 .power_up = "low";

dffeas \mem~145 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~145_q ),
	.prn(vcc));
defparam \mem~145 .is_wysiwyg = "true";
defparam \mem~145 .power_up = "low";

cycloneive_lcell_comb \mem~381 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~209_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~145_q ),
	.cin(gnd),
	.combout(\mem~381_combout ),
	.cout());
defparam \mem~381 .lut_mask = 16'hFFDE;
defparam \mem~381 .sum_lutc_input = "datac";

dffeas \mem~241 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~241_q ),
	.prn(vcc));
defparam \mem~241 .is_wysiwyg = "true";
defparam \mem~241 .power_up = "low";

cycloneive_lcell_comb \mem~382 (
	.dataa(\mem~177_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~381_combout ),
	.datad(\mem~241_q ),
	.cin(gnd),
	.combout(\mem~382_combout ),
	.cout());
defparam \mem~382 .lut_mask = 16'hFFBE;
defparam \mem~382 .sum_lutc_input = "datac";

dffeas \mem~81 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~81_q ),
	.prn(vcc));
defparam \mem~81 .is_wysiwyg = "true";
defparam \mem~81 .power_up = "low";

dffeas \mem~49 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~49_q ),
	.prn(vcc));
defparam \mem~49 .is_wysiwyg = "true";
defparam \mem~49 .power_up = "low";

dffeas \mem~17 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~17_q ),
	.prn(vcc));
defparam \mem~17 .is_wysiwyg = "true";
defparam \mem~17 .power_up = "low";

cycloneive_lcell_comb \mem~383 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~49_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~17_q ),
	.cin(gnd),
	.combout(\mem~383_combout ),
	.cout());
defparam \mem~383 .lut_mask = 16'hFFDE;
defparam \mem~383 .sum_lutc_input = "datac";

dffeas \mem~113 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~113_q ),
	.prn(vcc));
defparam \mem~113 .is_wysiwyg = "true";
defparam \mem~113 .power_up = "low";

cycloneive_lcell_comb \mem~384 (
	.dataa(\mem~81_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~383_combout ),
	.datad(\mem~113_q ),
	.cin(gnd),
	.combout(\mem~384_combout ),
	.cout());
defparam \mem~384 .lut_mask = 16'hFFBE;
defparam \mem~384 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~385 (
	.dataa(\mem~382_combout ),
	.datab(\mem~384_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~385_combout ),
	.cout());
defparam \mem~385 .lut_mask = 16'hAACC;
defparam \mem~385 .sum_lutc_input = "datac";

dffeas \internal_out_payload[17] (
	.clk(clk),
	.d(\mem~385_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[17]~q ),
	.prn(vcc));
defparam \internal_out_payload[17] .is_wysiwyg = "true";
defparam \internal_out_payload[17] .power_up = "low";

dffeas \mem~181 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~181_q ),
	.prn(vcc));
defparam \mem~181 .is_wysiwyg = "true";
defparam \mem~181 .power_up = "low";

dffeas \mem~213 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~213_q ),
	.prn(vcc));
defparam \mem~213 .is_wysiwyg = "true";
defparam \mem~213 .power_up = "low";

dffeas \mem~149 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~149_q ),
	.prn(vcc));
defparam \mem~149 .is_wysiwyg = "true";
defparam \mem~149 .power_up = "low";

cycloneive_lcell_comb \mem~386 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~213_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~149_q ),
	.cin(gnd),
	.combout(\mem~386_combout ),
	.cout());
defparam \mem~386 .lut_mask = 16'hFFDE;
defparam \mem~386 .sum_lutc_input = "datac";

dffeas \mem~245 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~245_q ),
	.prn(vcc));
defparam \mem~245 .is_wysiwyg = "true";
defparam \mem~245 .power_up = "low";

cycloneive_lcell_comb \mem~387 (
	.dataa(\mem~181_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~386_combout ),
	.datad(\mem~245_q ),
	.cin(gnd),
	.combout(\mem~387_combout ),
	.cout());
defparam \mem~387 .lut_mask = 16'hFFBE;
defparam \mem~387 .sum_lutc_input = "datac";

dffeas \mem~85 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~85_q ),
	.prn(vcc));
defparam \mem~85 .is_wysiwyg = "true";
defparam \mem~85 .power_up = "low";

dffeas \mem~53 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~53_q ),
	.prn(vcc));
defparam \mem~53 .is_wysiwyg = "true";
defparam \mem~53 .power_up = "low";

dffeas \mem~21 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~21_q ),
	.prn(vcc));
defparam \mem~21 .is_wysiwyg = "true";
defparam \mem~21 .power_up = "low";

cycloneive_lcell_comb \mem~388 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~53_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~21_q ),
	.cin(gnd),
	.combout(\mem~388_combout ),
	.cout());
defparam \mem~388 .lut_mask = 16'hFFDE;
defparam \mem~388 .sum_lutc_input = "datac";

dffeas \mem~117 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~117_q ),
	.prn(vcc));
defparam \mem~117 .is_wysiwyg = "true";
defparam \mem~117 .power_up = "low";

cycloneive_lcell_comb \mem~389 (
	.dataa(\mem~85_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~388_combout ),
	.datad(\mem~117_q ),
	.cin(gnd),
	.combout(\mem~389_combout ),
	.cout());
defparam \mem~389 .lut_mask = 16'hFFBE;
defparam \mem~389 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~390 (
	.dataa(\mem~387_combout ),
	.datab(\mem~389_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~390_combout ),
	.cout());
defparam \mem~390 .lut_mask = 16'hAACC;
defparam \mem~390 .sum_lutc_input = "datac";

dffeas \internal_out_payload[21] (
	.clk(clk),
	.d(\mem~390_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[21]~q ),
	.prn(vcc));
defparam \internal_out_payload[21] .is_wysiwyg = "true";
defparam \internal_out_payload[21] .power_up = "low";

dffeas \mem~187 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~187_q ),
	.prn(vcc));
defparam \mem~187 .is_wysiwyg = "true";
defparam \mem~187 .power_up = "low";

dffeas \mem~219 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~219_q ),
	.prn(vcc));
defparam \mem~219 .is_wysiwyg = "true";
defparam \mem~219 .power_up = "low";

dffeas \mem~155 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~155_q ),
	.prn(vcc));
defparam \mem~155 .is_wysiwyg = "true";
defparam \mem~155 .power_up = "low";

cycloneive_lcell_comb \mem~391 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~219_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~155_q ),
	.cin(gnd),
	.combout(\mem~391_combout ),
	.cout());
defparam \mem~391 .lut_mask = 16'hFFDE;
defparam \mem~391 .sum_lutc_input = "datac";

dffeas \mem~251 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~251_q ),
	.prn(vcc));
defparam \mem~251 .is_wysiwyg = "true";
defparam \mem~251 .power_up = "low";

cycloneive_lcell_comb \mem~392 (
	.dataa(\mem~187_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~391_combout ),
	.datad(\mem~251_q ),
	.cin(gnd),
	.combout(\mem~392_combout ),
	.cout());
defparam \mem~392 .lut_mask = 16'hFFBE;
defparam \mem~392 .sum_lutc_input = "datac";

dffeas \mem~91 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~91_q ),
	.prn(vcc));
defparam \mem~91 .is_wysiwyg = "true";
defparam \mem~91 .power_up = "low";

dffeas \mem~59 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~59_q ),
	.prn(vcc));
defparam \mem~59 .is_wysiwyg = "true";
defparam \mem~59 .power_up = "low";

dffeas \mem~27 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~27_q ),
	.prn(vcc));
defparam \mem~27 .is_wysiwyg = "true";
defparam \mem~27 .power_up = "low";

cycloneive_lcell_comb \mem~393 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~59_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~27_q ),
	.cin(gnd),
	.combout(\mem~393_combout ),
	.cout());
defparam \mem~393 .lut_mask = 16'hFFDE;
defparam \mem~393 .sum_lutc_input = "datac";

dffeas \mem~123 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~123_q ),
	.prn(vcc));
defparam \mem~123 .is_wysiwyg = "true";
defparam \mem~123 .power_up = "low";

cycloneive_lcell_comb \mem~394 (
	.dataa(\mem~91_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~393_combout ),
	.datad(\mem~123_q ),
	.cin(gnd),
	.combout(\mem~394_combout ),
	.cout());
defparam \mem~394 .lut_mask = 16'hFFBE;
defparam \mem~394 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~395 (
	.dataa(\mem~392_combout ),
	.datab(\mem~394_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~395_combout ),
	.cout());
defparam \mem~395 .lut_mask = 16'hAACC;
defparam \mem~395 .sum_lutc_input = "datac";

dffeas \internal_out_payload[27] (
	.clk(clk),
	.d(\mem~395_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[27]~q ),
	.prn(vcc));
defparam \internal_out_payload[27] .is_wysiwyg = "true";
defparam \internal_out_payload[27] .power_up = "low";

dffeas \mem~188 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~188_q ),
	.prn(vcc));
defparam \mem~188 .is_wysiwyg = "true";
defparam \mem~188 .power_up = "low";

dffeas \mem~220 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~220_q ),
	.prn(vcc));
defparam \mem~220 .is_wysiwyg = "true";
defparam \mem~220 .power_up = "low";

dffeas \mem~156 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~156_q ),
	.prn(vcc));
defparam \mem~156 .is_wysiwyg = "true";
defparam \mem~156 .power_up = "low";

cycloneive_lcell_comb \mem~396 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~220_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~156_q ),
	.cin(gnd),
	.combout(\mem~396_combout ),
	.cout());
defparam \mem~396 .lut_mask = 16'hFFDE;
defparam \mem~396 .sum_lutc_input = "datac";

dffeas \mem~252 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~252_q ),
	.prn(vcc));
defparam \mem~252 .is_wysiwyg = "true";
defparam \mem~252 .power_up = "low";

cycloneive_lcell_comb \mem~397 (
	.dataa(\mem~188_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~396_combout ),
	.datad(\mem~252_q ),
	.cin(gnd),
	.combout(\mem~397_combout ),
	.cout());
defparam \mem~397 .lut_mask = 16'hFFBE;
defparam \mem~397 .sum_lutc_input = "datac";

dffeas \mem~92 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~92_q ),
	.prn(vcc));
defparam \mem~92 .is_wysiwyg = "true";
defparam \mem~92 .power_up = "low";

dffeas \mem~60 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~60_q ),
	.prn(vcc));
defparam \mem~60 .is_wysiwyg = "true";
defparam \mem~60 .power_up = "low";

dffeas \mem~28 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~28_q ),
	.prn(vcc));
defparam \mem~28 .is_wysiwyg = "true";
defparam \mem~28 .power_up = "low";

cycloneive_lcell_comb \mem~398 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~60_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~28_q ),
	.cin(gnd),
	.combout(\mem~398_combout ),
	.cout());
defparam \mem~398 .lut_mask = 16'hFFDE;
defparam \mem~398 .sum_lutc_input = "datac";

dffeas \mem~124 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~124_q ),
	.prn(vcc));
defparam \mem~124 .is_wysiwyg = "true";
defparam \mem~124 .power_up = "low";

cycloneive_lcell_comb \mem~399 (
	.dataa(\mem~92_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~398_combout ),
	.datad(\mem~124_q ),
	.cin(gnd),
	.combout(\mem~399_combout ),
	.cout());
defparam \mem~399 .lut_mask = 16'hFFBE;
defparam \mem~399 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~400 (
	.dataa(\mem~397_combout ),
	.datab(\mem~399_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~400_combout ),
	.cout());
defparam \mem~400 .lut_mask = 16'hAACC;
defparam \mem~400 .sum_lutc_input = "datac";

dffeas \internal_out_payload[28] (
	.clk(clk),
	.d(\mem~400_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[28]~q ),
	.prn(vcc));
defparam \internal_out_payload[28] .is_wysiwyg = "true";
defparam \internal_out_payload[28] .power_up = "low";

dffeas \mem~191 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~191_q ),
	.prn(vcc));
defparam \mem~191 .is_wysiwyg = "true";
defparam \mem~191 .power_up = "low";

dffeas \mem~223 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~223_q ),
	.prn(vcc));
defparam \mem~223 .is_wysiwyg = "true";
defparam \mem~223 .power_up = "low";

dffeas \mem~159 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~159_q ),
	.prn(vcc));
defparam \mem~159 .is_wysiwyg = "true";
defparam \mem~159 .power_up = "low";

cycloneive_lcell_comb \mem~401 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~223_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~159_q ),
	.cin(gnd),
	.combout(\mem~401_combout ),
	.cout());
defparam \mem~401 .lut_mask = 16'hFFDE;
defparam \mem~401 .sum_lutc_input = "datac";

dffeas \mem~255 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~255_q ),
	.prn(vcc));
defparam \mem~255 .is_wysiwyg = "true";
defparam \mem~255 .power_up = "low";

cycloneive_lcell_comb \mem~402 (
	.dataa(\mem~191_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~401_combout ),
	.datad(\mem~255_q ),
	.cin(gnd),
	.combout(\mem~402_combout ),
	.cout());
defparam \mem~402 .lut_mask = 16'hFFBE;
defparam \mem~402 .sum_lutc_input = "datac";

dffeas \mem~95 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~95_q ),
	.prn(vcc));
defparam \mem~95 .is_wysiwyg = "true";
defparam \mem~95 .power_up = "low";

dffeas \mem~63 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~63_q ),
	.prn(vcc));
defparam \mem~63 .is_wysiwyg = "true";
defparam \mem~63 .power_up = "low";

dffeas \mem~31 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~31_q ),
	.prn(vcc));
defparam \mem~31 .is_wysiwyg = "true";
defparam \mem~31 .power_up = "low";

cycloneive_lcell_comb \mem~403 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~63_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~31_q ),
	.cin(gnd),
	.combout(\mem~403_combout ),
	.cout());
defparam \mem~403 .lut_mask = 16'hFFDE;
defparam \mem~403 .sum_lutc_input = "datac";

dffeas \mem~127 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~127_q ),
	.prn(vcc));
defparam \mem~127 .is_wysiwyg = "true";
defparam \mem~127 .power_up = "low";

cycloneive_lcell_comb \mem~404 (
	.dataa(\mem~95_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~403_combout ),
	.datad(\mem~127_q ),
	.cin(gnd),
	.combout(\mem~404_combout ),
	.cout());
defparam \mem~404 .lut_mask = 16'hFFBE;
defparam \mem~404 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~405 (
	.dataa(\mem~402_combout ),
	.datab(\mem~404_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~405_combout ),
	.cout());
defparam \mem~405 .lut_mask = 16'hAACC;
defparam \mem~405 .sum_lutc_input = "datac";

dffeas \internal_out_payload[31] (
	.clk(clk),
	.d(\mem~405_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[31]~q ),
	.prn(vcc));
defparam \internal_out_payload[31] .is_wysiwyg = "true";
defparam \internal_out_payload[31] .power_up = "low";

dffeas \mem~190 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~190_q ),
	.prn(vcc));
defparam \mem~190 .is_wysiwyg = "true";
defparam \mem~190 .power_up = "low";

dffeas \mem~222 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~222_q ),
	.prn(vcc));
defparam \mem~222 .is_wysiwyg = "true";
defparam \mem~222 .power_up = "low";

dffeas \mem~158 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~158_q ),
	.prn(vcc));
defparam \mem~158 .is_wysiwyg = "true";
defparam \mem~158 .power_up = "low";

cycloneive_lcell_comb \mem~406 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~222_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~158_q ),
	.cin(gnd),
	.combout(\mem~406_combout ),
	.cout());
defparam \mem~406 .lut_mask = 16'hFFDE;
defparam \mem~406 .sum_lutc_input = "datac";

dffeas \mem~254 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~254_q ),
	.prn(vcc));
defparam \mem~254 .is_wysiwyg = "true";
defparam \mem~254 .power_up = "low";

cycloneive_lcell_comb \mem~407 (
	.dataa(\mem~190_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~406_combout ),
	.datad(\mem~254_q ),
	.cin(gnd),
	.combout(\mem~407_combout ),
	.cout());
defparam \mem~407 .lut_mask = 16'hFFBE;
defparam \mem~407 .sum_lutc_input = "datac";

dffeas \mem~94 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~94_q ),
	.prn(vcc));
defparam \mem~94 .is_wysiwyg = "true";
defparam \mem~94 .power_up = "low";

dffeas \mem~62 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~62_q ),
	.prn(vcc));
defparam \mem~62 .is_wysiwyg = "true";
defparam \mem~62 .power_up = "low";

dffeas \mem~30 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~30_q ),
	.prn(vcc));
defparam \mem~30 .is_wysiwyg = "true";
defparam \mem~30 .power_up = "low";

cycloneive_lcell_comb \mem~408 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~62_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~30_q ),
	.cin(gnd),
	.combout(\mem~408_combout ),
	.cout());
defparam \mem~408 .lut_mask = 16'hFFDE;
defparam \mem~408 .sum_lutc_input = "datac";

dffeas \mem~126 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~126_q ),
	.prn(vcc));
defparam \mem~126 .is_wysiwyg = "true";
defparam \mem~126 .power_up = "low";

cycloneive_lcell_comb \mem~409 (
	.dataa(\mem~94_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~408_combout ),
	.datad(\mem~126_q ),
	.cin(gnd),
	.combout(\mem~409_combout ),
	.cout());
defparam \mem~409 .lut_mask = 16'hFFBE;
defparam \mem~409 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~410 (
	.dataa(\mem~407_combout ),
	.datab(\mem~409_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~410_combout ),
	.cout());
defparam \mem~410 .lut_mask = 16'hAACC;
defparam \mem~410 .sum_lutc_input = "datac";

dffeas \internal_out_payload[30] (
	.clk(clk),
	.d(\mem~410_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[30]~q ),
	.prn(vcc));
defparam \internal_out_payload[30] .is_wysiwyg = "true";
defparam \internal_out_payload[30] .power_up = "low";

dffeas \mem~189 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~189_q ),
	.prn(vcc));
defparam \mem~189 .is_wysiwyg = "true";
defparam \mem~189 .power_up = "low";

dffeas \mem~221 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~221_q ),
	.prn(vcc));
defparam \mem~221 .is_wysiwyg = "true";
defparam \mem~221 .power_up = "low";

dffeas \mem~157 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~157_q ),
	.prn(vcc));
defparam \mem~157 .is_wysiwyg = "true";
defparam \mem~157 .power_up = "low";

cycloneive_lcell_comb \mem~411 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~221_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~157_q ),
	.cin(gnd),
	.combout(\mem~411_combout ),
	.cout());
defparam \mem~411 .lut_mask = 16'hFFDE;
defparam \mem~411 .sum_lutc_input = "datac";

dffeas \mem~253 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~253_q ),
	.prn(vcc));
defparam \mem~253 .is_wysiwyg = "true";
defparam \mem~253 .power_up = "low";

cycloneive_lcell_comb \mem~412 (
	.dataa(\mem~189_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~411_combout ),
	.datad(\mem~253_q ),
	.cin(gnd),
	.combout(\mem~412_combout ),
	.cout());
defparam \mem~412 .lut_mask = 16'hFFBE;
defparam \mem~412 .sum_lutc_input = "datac";

dffeas \mem~93 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~93_q ),
	.prn(vcc));
defparam \mem~93 .is_wysiwyg = "true";
defparam \mem~93 .power_up = "low";

dffeas \mem~61 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~61_q ),
	.prn(vcc));
defparam \mem~61 .is_wysiwyg = "true";
defparam \mem~61 .power_up = "low";

dffeas \mem~29 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~29_q ),
	.prn(vcc));
defparam \mem~29 .is_wysiwyg = "true";
defparam \mem~29 .power_up = "low";

cycloneive_lcell_comb \mem~413 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~61_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~29_q ),
	.cin(gnd),
	.combout(\mem~413_combout ),
	.cout());
defparam \mem~413 .lut_mask = 16'hFFDE;
defparam \mem~413 .sum_lutc_input = "datac";

dffeas \mem~125 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~125_q ),
	.prn(vcc));
defparam \mem~125 .is_wysiwyg = "true";
defparam \mem~125 .power_up = "low";

cycloneive_lcell_comb \mem~414 (
	.dataa(\mem~93_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~413_combout ),
	.datad(\mem~125_q ),
	.cin(gnd),
	.combout(\mem~414_combout ),
	.cout());
defparam \mem~414 .lut_mask = 16'hFFBE;
defparam \mem~414 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~415 (
	.dataa(\mem~412_combout ),
	.datab(\mem~414_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~415_combout ),
	.cout());
defparam \mem~415 .lut_mask = 16'hAACC;
defparam \mem~415 .sum_lutc_input = "datac";

dffeas \internal_out_payload[29] (
	.clk(clk),
	.d(\mem~415_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[29]~q ),
	.prn(vcc));
defparam \internal_out_payload[29] .is_wysiwyg = "true";
defparam \internal_out_payload[29] .power_up = "low";

endmodule

module usb_system_altera_avalon_sc_fifo_9 (
	clk,
	reset,
	mem_used_7,
	last_cycle,
	saved_grant_0,
	saved_grant_1,
	WideOr1,
	out_data_buffer_67,
	src_data_68,
	nonposted_write_endofpacket,
	mem_used_0,
	mem_107_0,
	out_valid,
	mem_86_0,
	mem_68_0,
	WideOr0,
	mem_67_0,
	out_data_buffer_86)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
output 	mem_used_7;
input 	last_cycle;
input 	saved_grant_0;
input 	saved_grant_1;
input 	WideOr1;
input 	out_data_buffer_67;
input 	src_data_68;
input 	nonposted_write_endofpacket;
output 	mem_used_0;
output 	mem_107_0;
input 	out_valid;
output 	mem_86_0;
output 	mem_68_0;
input 	WideOr0;
output 	mem_67_0;
input 	out_data_buffer_86;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used~6_combout ;
wire \read~0_combout ;
wire \mem_used[6]~2_combout ;
wire \mem_used[1]~q ;
wire \mem_used~8_combout ;
wire \mem_used[2]~q ;
wire \mem_used~9_combout ;
wire \mem_used[3]~q ;
wire \mem_used~7_combout ;
wire \mem_used[4]~q ;
wire \mem_used~5_combout ;
wire \mem_used[5]~q ;
wire \mem_used~1_combout ;
wire \mem_used[6]~q ;
wire \mem_used[7]~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem[7][107]~q ;
wire \mem~24_combout ;
wire \always6~0_combout ;
wire \mem[6][107]~q ;
wire \mem~20_combout ;
wire \always5~0_combout ;
wire \mem[5][107]~q ;
wire \mem~16_combout ;
wire \always4~0_combout ;
wire \mem[4][107]~q ;
wire \mem~12_combout ;
wire \always3~0_combout ;
wire \mem[3][107]~q ;
wire \mem~8_combout ;
wire \always2~0_combout ;
wire \mem[2][107]~q ;
wire \mem~4_combout ;
wire \always1~0_combout ;
wire \mem[1][107]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[7][86]~q ;
wire \mem~25_combout ;
wire \mem[6][86]~q ;
wire \mem~21_combout ;
wire \mem[5][86]~q ;
wire \mem~17_combout ;
wire \mem[4][86]~q ;
wire \mem~13_combout ;
wire \mem[3][86]~q ;
wire \mem~9_combout ;
wire \mem[2][86]~q ;
wire \mem~5_combout ;
wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem[7][68]~q ;
wire \mem~26_combout ;
wire \mem[6][68]~q ;
wire \mem~22_combout ;
wire \mem[5][68]~q ;
wire \mem~18_combout ;
wire \mem[4][68]~q ;
wire \mem~14_combout ;
wire \mem[3][68]~q ;
wire \mem~10_combout ;
wire \mem[2][68]~q ;
wire \mem~6_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;
wire \mem[7][67]~q ;
wire \mem~27_combout ;
wire \mem[6][67]~q ;
wire \mem~23_combout ;
wire \mem[5][67]~q ;
wire \mem~19_combout ;
wire \mem[4][67]~q ;
wire \mem~15_combout ;
wire \mem[3][67]~q ;
wire \mem~11_combout ;
wire \mem[2][67]~q ;
wire \mem~7_combout ;
wire \mem[1][67]~q ;
wire \mem~3_combout ;


dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used[7]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_7),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(last_cycle),
	.datab(nonposted_write_endofpacket),
	.datac(WideOr1),
	.datad(src_data_68),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFFFE;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used~6 (
	.dataa(mem_used_0),
	.datab(\mem_used[2]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~6_combout ),
	.cout());
defparam \mem_used~6 .lut_mask = 16'hAACC;
defparam \mem_used~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(mem_used_0),
	.datab(mem_107_0),
	.datac(out_valid),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hFEFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[6]~2 (
	.dataa(\write~0_combout ),
	.datab(\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[6]~2_combout ),
	.cout());
defparam \mem_used[6]~2 .lut_mask = 16'h6666;
defparam \mem_used[6]~2 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used~8 (
	.dataa(\mem_used[1]~q ),
	.datab(\mem_used[3]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~8_combout ),
	.cout());
defparam \mem_used~8 .lut_mask = 16'hAACC;
defparam \mem_used~8 .sum_lutc_input = "datac";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cycloneive_lcell_comb \mem_used~9 (
	.dataa(\mem_used[2]~q ),
	.datab(\mem_used[4]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~9_combout ),
	.cout());
defparam \mem_used~9 .lut_mask = 16'hAACC;
defparam \mem_used~9 .sum_lutc_input = "datac";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cycloneive_lcell_comb \mem_used~7 (
	.dataa(\mem_used[3]~q ),
	.datab(\mem_used[5]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~7_combout ),
	.cout());
defparam \mem_used~7 .lut_mask = 16'hAACC;
defparam \mem_used~7 .sum_lutc_input = "datac";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cycloneive_lcell_comb \mem_used~5 (
	.dataa(\mem_used[4]~q ),
	.datab(\mem_used[6]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~5_combout ),
	.cout());
defparam \mem_used~5 .lut_mask = 16'hAACC;
defparam \mem_used~5 .sum_lutc_input = "datac";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cycloneive_lcell_comb \mem_used~1 (
	.dataa(mem_used_7),
	.datab(\write~0_combout ),
	.datac(\mem_used[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used~1_combout ),
	.cout());
defparam \mem_used~1 .lut_mask = 16'hFEFE;
defparam \mem_used~1 .sum_lutc_input = "datac";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cycloneive_lcell_comb \mem_used[7]~0 (
	.dataa(mem_used_7),
	.datab(\write~0_combout ),
	.datac(\mem_used[6]~q ),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[7]~0_combout ),
	.cout());
defparam \mem_used[7]~0 .lut_mask = 16'hFBFE;
defparam \mem_used[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[1]~q ),
	.datab(gnd),
	.datac(mem_107_0),
	.datad(out_valid),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hAFFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\write~0_combout ),
	.datab(mem_used_0),
	.datac(WideOr0),
	.datad(\mem_used[0]~3_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem[7][107] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][107]~q ),
	.prn(vcc));
defparam \mem[7][107] .is_wysiwyg = "true";
defparam \mem[7][107] .power_up = "low";

cycloneive_lcell_comb \mem~24 (
	.dataa(\mem[7][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~24_combout ),
	.cout());
defparam \mem~24 .lut_mask = 16'hAACC;
defparam \mem~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always6~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\always6~0_combout ),
	.cout());
defparam \always6~0 .lut_mask = 16'hAAFF;
defparam \always6~0 .sum_lutc_input = "datac";

dffeas \mem[6][107] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][107]~q ),
	.prn(vcc));
defparam \mem[6][107] .is_wysiwyg = "true";
defparam \mem[6][107] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[6][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'hAAFF;
defparam \always5~0 .sum_lutc_input = "datac";

dffeas \mem[5][107] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][107]~q ),
	.prn(vcc));
defparam \mem[5][107] .is_wysiwyg = "true";
defparam \mem[5][107] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[5][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAACC;
defparam \mem~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hAAFF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas \mem[4][107] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][107]~q ),
	.prn(vcc));
defparam \mem[4][107] .is_wysiwyg = "true";
defparam \mem[4][107] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[4][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always3~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hAAFF;
defparam \always3~0 .sum_lutc_input = "datac";

dffeas \mem[3][107] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][107]~q ),
	.prn(vcc));
defparam \mem[3][107] .is_wysiwyg = "true";
defparam \mem[3][107] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[3][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hAACC;
defparam \mem~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

dffeas \mem[2][107] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][107]~q ),
	.prn(vcc));
defparam \mem[2][107] .is_wysiwyg = "true";
defparam \mem[2][107] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[2][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hAAFF;
defparam \always1~0 .sum_lutc_input = "datac";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(mem_107_0),
	.datab(out_valid),
	.datac(WideOr0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hEFFF;
defparam \always0~0 .sum_lutc_input = "datac";

dffeas \mem[7][86] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][86]~q ),
	.prn(vcc));
defparam \mem[7][86] .is_wysiwyg = "true";
defparam \mem[7][86] .power_up = "low";

cycloneive_lcell_comb \mem~25 (
	.dataa(\mem[7][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~25_combout ),
	.cout());
defparam \mem~25 .lut_mask = 16'hFAFC;
defparam \mem~25 .sum_lutc_input = "datac";

dffeas \mem[6][86] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][86]~q ),
	.prn(vcc));
defparam \mem[6][86] .is_wysiwyg = "true";
defparam \mem[6][86] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[6][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hFAFC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[5][86] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][86]~q ),
	.prn(vcc));
defparam \mem[5][86] .is_wysiwyg = "true";
defparam \mem[5][86] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[5][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hFAFC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[4][86] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][86]~q ),
	.prn(vcc));
defparam \mem[4][86] .is_wysiwyg = "true";
defparam \mem[4][86] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[4][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hFAFC;
defparam \mem~13 .sum_lutc_input = "datac";

dffeas \mem[3][86] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][86]~q ),
	.prn(vcc));
defparam \mem[3][86] .is_wysiwyg = "true";
defparam \mem[3][86] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[3][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hFAFC;
defparam \mem~9 .sum_lutc_input = "datac";

dffeas \mem[2][86] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][86]~q ),
	.prn(vcc));
defparam \mem[2][86] .is_wysiwyg = "true";
defparam \mem[2][86] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[2][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hFAFC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hFAFC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[7][68] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][68]~q ),
	.prn(vcc));
defparam \mem[7][68] .is_wysiwyg = "true";
defparam \mem[7][68] .power_up = "low";

cycloneive_lcell_comb \mem~26 (
	.dataa(\mem[7][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~26_combout ),
	.cout());
defparam \mem~26 .lut_mask = 16'hAACC;
defparam \mem~26 .sum_lutc_input = "datac";

dffeas \mem[6][68] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][68]~q ),
	.prn(vcc));
defparam \mem[6][68] .is_wysiwyg = "true";
defparam \mem[6][68] .power_up = "low";

cycloneive_lcell_comb \mem~22 (
	.dataa(\mem[6][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~22_combout ),
	.cout());
defparam \mem~22 .lut_mask = 16'hAACC;
defparam \mem~22 .sum_lutc_input = "datac";

dffeas \mem[5][68] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][68]~q ),
	.prn(vcc));
defparam \mem[5][68] .is_wysiwyg = "true";
defparam \mem[5][68] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[5][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

dffeas \mem[4][68] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][68]~q ),
	.prn(vcc));
defparam \mem[4][68] .is_wysiwyg = "true";
defparam \mem[4][68] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[4][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[3][68] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][68]~q ),
	.prn(vcc));
defparam \mem[3][68] .is_wysiwyg = "true";
defparam \mem[3][68] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[3][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hAACC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[2][68] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][68]~q ),
	.prn(vcc));
defparam \mem[2][68] .is_wysiwyg = "true";
defparam \mem[2][68] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[2][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[7][67] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][67]~q ),
	.prn(vcc));
defparam \mem[7][67] .is_wysiwyg = "true";
defparam \mem[7][67] .power_up = "low";

cycloneive_lcell_comb \mem~27 (
	.dataa(\mem[7][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~27_combout ),
	.cout());
defparam \mem~27 .lut_mask = 16'hFAFC;
defparam \mem~27 .sum_lutc_input = "datac";

dffeas \mem[6][67] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][67]~q ),
	.prn(vcc));
defparam \mem[6][67] .is_wysiwyg = "true";
defparam \mem[6][67] .power_up = "low";

cycloneive_lcell_comb \mem~23 (
	.dataa(\mem[6][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~23_combout ),
	.cout());
defparam \mem~23 .lut_mask = 16'hFAFC;
defparam \mem~23 .sum_lutc_input = "datac";

dffeas \mem[5][67] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][67]~q ),
	.prn(vcc));
defparam \mem[5][67] .is_wysiwyg = "true";
defparam \mem[5][67] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[5][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hFAFC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[4][67] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][67]~q ),
	.prn(vcc));
defparam \mem[4][67] .is_wysiwyg = "true";
defparam \mem[4][67] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[4][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hFAFC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[3][67] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][67]~q ),
	.prn(vcc));
defparam \mem[3][67] .is_wysiwyg = "true";
defparam \mem[3][67] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[3][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hFAFC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[2][67] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][67]~q ),
	.prn(vcc));
defparam \mem[2][67] .is_wysiwyg = "true";
defparam \mem[2][67] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[2][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hFAFC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFAFC;
defparam \mem~3 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_sc_fifo_10 (
	reset,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	uav_write,
	saved_grant_0,
	saved_grant_1,
	mem_used_1,
	src_data_68,
	read_latency_shift_reg,
	WideOr1,
	cp_ready,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	uav_write;
input 	saved_grant_0;
input 	saved_grant_1;
output 	mem_used_1;
input 	src_data_68;
input 	read_latency_shift_reg;
input 	WideOr1;
input 	cp_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~1_combout ;
wire \mem[1][67]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~2_combout ),
	.datab(WideOr1),
	.datac(src_data_68),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hFAFC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hACFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_avalon_st_handshake_clock_crosser (
	wire_pll7_clk_0,
	W_alu_result_7,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_8,
	W_alu_result_6,
	W_alu_result_24,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	altera_reset_synchronizer_int_chain_out,
	uav_write,
	uav_read,
	sink_ready,
	in_data_toggle,
	dreg_0,
	s0_cmd_valid,
	last_cycle,
	saved_grant_0,
	out_data_toggle_flopped,
	dreg_01,
	out_valid,
	out_data_buffer_67,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	sink_ready1,
	out_data_buffer_107,
	out_data_buffer_66,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_18,
	out_data_buffer_19,
	out_data_buffer_20,
	out_data_buffer_21,
	out_data_buffer_22,
	out_data_buffer_23,
	out_data_buffer_24,
	out_data_buffer_25,
	out_data_buffer_26,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_29,
	out_data_buffer_30,
	out_data_buffer_31,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_7;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_8;
input 	W_alu_result_6;
input 	W_alu_result_24;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	altera_reset_synchronizer_int_chain_out;
input 	uav_write;
input 	uav_read;
input 	sink_ready;
output 	in_data_toggle;
output 	dreg_0;
input 	s0_cmd_valid;
input 	last_cycle;
input 	saved_grant_0;
output 	out_data_toggle_flopped;
output 	dreg_01;
output 	out_valid;
output 	out_data_buffer_67;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
input 	sink_ready1;
output 	out_data_buffer_107;
output 	out_data_buffer_66;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_18;
output 	out_data_buffer_19;
output 	out_data_buffer_20;
output 	out_data_buffer_21;
output 	out_data_buffer_22;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_29;
output 	out_data_buffer_30;
output 	out_data_buffer_31;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_avalon_st_clock_crosser_3 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,uav_write,uav_write,gnd,gnd,gnd,W_alu_result_26,W_alu_result_25,W_alu_result_24,W_alu_result_23,
W_alu_result_22,W_alu_result_21,W_alu_result_20,W_alu_result_19,W_alu_result_18,W_alu_result_17,W_alu_result_16,W_alu_result_15,W_alu_result_14,W_alu_result_13,W_alu_result_12,W_alu_result_11,W_alu_result_10,W_alu_result_9,W_alu_result_8,W_alu_result_7,W_alu_result_6,
W_alu_result_5,W_alu_result_4,W_alu_result_3,W_alu_result_2,gnd,gnd,d_byteenable_3,d_byteenable_2,d_byteenable_1,d_byteenable_0,d_writedata_31,d_writedata_30,d_writedata_29,d_writedata_28,d_writedata_27,d_writedata_26,d_writedata_25,d_writedata_24,d_writedata_23,
d_writedata_22,d_writedata_21,d_writedata_20,d_writedata_19,d_writedata_18,d_writedata_17,d_writedata_16,d_writedata_15,d_writedata_14,d_writedata_13,d_writedata_12,d_writedata_11,d_writedata_10,d_writedata_9,d_writedata_8,d_writedata_7,d_writedata_6,d_writedata_5,
d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.in_reset(r_sync_rst),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.sink_ready(sink_ready),
	.in_data_toggle1(in_data_toggle),
	.dreg_0(dreg_0),
	.s0_cmd_valid(s0_cmd_valid),
	.last_cycle(last_cycle),
	.saved_grant_0(saved_grant_0),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_01(dreg_01),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_68(out_data_buffer_68),
	.out_data_buffer_48(out_data_buffer_48),
	.out_data_buffer_62(out_data_buffer_62),
	.out_data_buffer_49(out_data_buffer_49),
	.out_data_buffer_51(out_data_buffer_51),
	.out_data_buffer_50(out_data_buffer_50),
	.out_data_buffer_53(out_data_buffer_53),
	.out_data_buffer_52(out_data_buffer_52),
	.out_data_buffer_55(out_data_buffer_55),
	.out_data_buffer_54(out_data_buffer_54),
	.out_data_buffer_57(out_data_buffer_57),
	.out_data_buffer_56(out_data_buffer_56),
	.out_data_buffer_59(out_data_buffer_59),
	.out_data_buffer_58(out_data_buffer_58),
	.out_data_buffer_61(out_data_buffer_61),
	.out_data_buffer_60(out_data_buffer_60),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_buffer_40(out_data_buffer_40),
	.out_data_buffer_41(out_data_buffer_41),
	.out_data_buffer_42(out_data_buffer_42),
	.out_data_buffer_43(out_data_buffer_43),
	.out_data_buffer_44(out_data_buffer_44),
	.out_data_buffer_45(out_data_buffer_45),
	.out_data_buffer_46(out_data_buffer_46),
	.out_data_buffer_47(out_data_buffer_47),
	.out_data_buffer_32(out_data_buffer_32),
	.out_data_buffer_33(out_data_buffer_33),
	.out_data_buffer_34(out_data_buffer_34),
	.out_data_buffer_35(out_data_buffer_35),
	.sink_ready1(sink_ready1),
	.out_data_buffer_107(out_data_buffer_107),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_31(out_data_buffer_31),
	.clk_clk(clk_clk));

endmodule

module usb_system_altera_avalon_st_handshake_clock_crosser_1 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_5,
	F_pc_6,
	F_pc_4,
	F_pc_1,
	F_pc_3,
	i_read,
	read_accepted,
	F_pc_2,
	Equal2,
	F_pc_0,
	last_cycle,
	saved_grant_1,
	out_valid,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	always1,
	Equal1,
	take_in_data,
	out_data_buffer_107,
	out_data_buffer_86,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_4;
input 	F_pc_1;
input 	F_pc_3;
input 	i_read;
input 	read_accepted;
input 	F_pc_2;
input 	Equal2;
input 	F_pc_0;
input 	last_cycle;
input 	saved_grant_1;
output 	out_valid;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
input 	always1;
input 	Equal1;
output 	take_in_data;
output 	out_data_buffer_107;
output 	out_data_buffer_86;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_avalon_st_clock_crosser clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_reset(r_sync_rst),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,F_pc_24,F_pc_23,F_pc_22,F_pc_21,F_pc_20,F_pc_19,F_pc_18,F_pc_17,F_pc_16,F_pc_15,F_pc_14,F_pc_13,
F_pc_12,F_pc_11,F_pc_10,F_pc_9,F_pc_8,F_pc_7,F_pc_6,F_pc_5,F_pc_4,F_pc_3,F_pc_2,F_pc_1,F_pc_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.i_read(i_read),
	.read_accepted(read_accepted),
	.Equal2(Equal2),
	.last_cycle(last_cycle),
	.saved_grant_1(saved_grant_1),
	.out_valid1(out_valid),
	.out_data_buffer_68(out_data_buffer_68),
	.out_data_buffer_48(out_data_buffer_48),
	.out_data_buffer_62(out_data_buffer_62),
	.out_data_buffer_49(out_data_buffer_49),
	.out_data_buffer_51(out_data_buffer_51),
	.out_data_buffer_50(out_data_buffer_50),
	.out_data_buffer_53(out_data_buffer_53),
	.out_data_buffer_52(out_data_buffer_52),
	.out_data_buffer_55(out_data_buffer_55),
	.out_data_buffer_54(out_data_buffer_54),
	.out_data_buffer_57(out_data_buffer_57),
	.out_data_buffer_56(out_data_buffer_56),
	.out_data_buffer_59(out_data_buffer_59),
	.out_data_buffer_58(out_data_buffer_58),
	.out_data_buffer_61(out_data_buffer_61),
	.out_data_buffer_60(out_data_buffer_60),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_buffer_40(out_data_buffer_40),
	.out_data_buffer_41(out_data_buffer_41),
	.out_data_buffer_42(out_data_buffer_42),
	.out_data_buffer_43(out_data_buffer_43),
	.out_data_buffer_44(out_data_buffer_44),
	.out_data_buffer_45(out_data_buffer_45),
	.out_data_buffer_46(out_data_buffer_46),
	.out_data_buffer_47(out_data_buffer_47),
	.out_data_buffer_32(out_data_buffer_32),
	.out_data_buffer_33(out_data_buffer_33),
	.out_data_buffer_34(out_data_buffer_34),
	.out_data_buffer_35(out_data_buffer_35),
	.always1(always1),
	.Equal1(Equal1),
	.take_in_data(take_in_data),
	.out_data_buffer_107(out_data_buffer_107),
	.out_data_buffer_86(out_data_buffer_86),
	.clk_clk(clk_clk));

endmodule

module usb_system_altera_avalon_st_clock_crosser (
	wire_pll7_clk_0,
	in_reset,
	out_reset,
	in_data,
	i_read,
	read_accepted,
	Equal2,
	last_cycle,
	saved_grant_1,
	out_valid1,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	always1,
	Equal1,
	take_in_data,
	out_data_buffer_107,
	out_data_buffer_86,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	in_reset;
input 	out_reset;
input 	[118:0] in_data;
input 	i_read;
input 	read_accepted;
input 	Equal2;
input 	last_cycle;
input 	saved_grant_1;
output 	out_valid1;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
input 	always1;
input 	Equal1;
output 	take_in_data;
output 	out_data_buffer_107;
output 	out_data_buffer_86;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_to_out_synchronizer|dreg[0]~q ;
wire \out_to_in_synchronizer|dreg[0]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \out_data_toggle_flopped~q ;
wire \take_in_data~3_combout ;
wire \in_data_buffer[68]~q ;
wire \in_data_buffer[48]~q ;
wire \in_data_buffer[62]~q ;
wire \in_data_buffer[49]~q ;
wire \in_data_buffer[51]~q ;
wire \in_data_buffer[50]~q ;
wire \in_data_buffer[53]~q ;
wire \in_data_buffer[52]~q ;
wire \in_data_buffer[55]~q ;
wire \in_data_buffer[54]~q ;
wire \in_data_buffer[57]~q ;
wire \in_data_buffer[56]~q ;
wire \in_data_buffer[59]~q ;
wire \in_data_buffer[58]~q ;
wire \in_data_buffer[61]~q ;
wire \in_data_buffer[60]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[40]~q ;
wire \in_data_buffer[41]~q ;
wire \in_data_buffer[42]~q ;
wire \in_data_buffer[43]~q ;
wire \in_data_buffer[44]~q ;
wire \in_data_buffer[45]~q ;
wire \in_data_buffer[46]~q ;
wire \in_data_buffer[47]~q ;
wire \in_data_buffer[32]~q ;
wire \in_data_buffer[33]~q ;
wire \in_data_buffer[34]~q ;
wire \in_data_buffer[35]~q ;
wire \in_data_toggle~2_combout ;
wire \in_data_toggle~q ;
wire \in_ready~0_combout ;
wire \in_data_buffer[107]~q ;
wire \in_data_buffer[86]~q ;


usb_system_altera_std_synchronizer_7 out_to_in_synchronizer(
	.reset_n(in_reset),
	.din(\out_data_toggle_flopped~q ),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_6 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.dreg_0(\in_to_out_synchronizer|dreg[0]~q ),
	.din(\in_data_toggle~q ));

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_data_toggle_flopped~q ),
	.datad(\in_to_out_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[68] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[68]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_68),
	.prn(vcc));
defparam \out_data_buffer[68] .is_wysiwyg = "true";
defparam \out_data_buffer[68] .power_up = "low";

dffeas \out_data_buffer[48] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[48]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_48),
	.prn(vcc));
defparam \out_data_buffer[48] .is_wysiwyg = "true";
defparam \out_data_buffer[48] .power_up = "low";

dffeas \out_data_buffer[62] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[62]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_62),
	.prn(vcc));
defparam \out_data_buffer[62] .is_wysiwyg = "true";
defparam \out_data_buffer[62] .power_up = "low";

dffeas \out_data_buffer[49] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[49]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_49),
	.prn(vcc));
defparam \out_data_buffer[49] .is_wysiwyg = "true";
defparam \out_data_buffer[49] .power_up = "low";

dffeas \out_data_buffer[51] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[51]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_51),
	.prn(vcc));
defparam \out_data_buffer[51] .is_wysiwyg = "true";
defparam \out_data_buffer[51] .power_up = "low";

dffeas \out_data_buffer[50] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[50]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_50),
	.prn(vcc));
defparam \out_data_buffer[50] .is_wysiwyg = "true";
defparam \out_data_buffer[50] .power_up = "low";

dffeas \out_data_buffer[53] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[53]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_53),
	.prn(vcc));
defparam \out_data_buffer[53] .is_wysiwyg = "true";
defparam \out_data_buffer[53] .power_up = "low";

dffeas \out_data_buffer[52] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[52]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_52),
	.prn(vcc));
defparam \out_data_buffer[52] .is_wysiwyg = "true";
defparam \out_data_buffer[52] .power_up = "low";

dffeas \out_data_buffer[55] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[55]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_55),
	.prn(vcc));
defparam \out_data_buffer[55] .is_wysiwyg = "true";
defparam \out_data_buffer[55] .power_up = "low";

dffeas \out_data_buffer[54] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[54]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_54),
	.prn(vcc));
defparam \out_data_buffer[54] .is_wysiwyg = "true";
defparam \out_data_buffer[54] .power_up = "low";

dffeas \out_data_buffer[57] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[57]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_57),
	.prn(vcc));
defparam \out_data_buffer[57] .is_wysiwyg = "true";
defparam \out_data_buffer[57] .power_up = "low";

dffeas \out_data_buffer[56] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[56]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_56),
	.prn(vcc));
defparam \out_data_buffer[56] .is_wysiwyg = "true";
defparam \out_data_buffer[56] .power_up = "low";

dffeas \out_data_buffer[59] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[59]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_59),
	.prn(vcc));
defparam \out_data_buffer[59] .is_wysiwyg = "true";
defparam \out_data_buffer[59] .power_up = "low";

dffeas \out_data_buffer[58] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[58]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_58),
	.prn(vcc));
defparam \out_data_buffer[58] .is_wysiwyg = "true";
defparam \out_data_buffer[58] .power_up = "low";

dffeas \out_data_buffer[61] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[61]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_61),
	.prn(vcc));
defparam \out_data_buffer[61] .is_wysiwyg = "true";
defparam \out_data_buffer[61] .power_up = "low";

dffeas \out_data_buffer[60] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[60]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_60),
	.prn(vcc));
defparam \out_data_buffer[60] .is_wysiwyg = "true";
defparam \out_data_buffer[60] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas \out_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[40]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_40),
	.prn(vcc));
defparam \out_data_buffer[40] .is_wysiwyg = "true";
defparam \out_data_buffer[40] .power_up = "low";

dffeas \out_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[41]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_41),
	.prn(vcc));
defparam \out_data_buffer[41] .is_wysiwyg = "true";
defparam \out_data_buffer[41] .power_up = "low";

dffeas \out_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[42]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_42),
	.prn(vcc));
defparam \out_data_buffer[42] .is_wysiwyg = "true";
defparam \out_data_buffer[42] .power_up = "low";

dffeas \out_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[43]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_43),
	.prn(vcc));
defparam \out_data_buffer[43] .is_wysiwyg = "true";
defparam \out_data_buffer[43] .power_up = "low";

dffeas \out_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[44]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_44),
	.prn(vcc));
defparam \out_data_buffer[44] .is_wysiwyg = "true";
defparam \out_data_buffer[44] .power_up = "low";

dffeas \out_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[45]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_45),
	.prn(vcc));
defparam \out_data_buffer[45] .is_wysiwyg = "true";
defparam \out_data_buffer[45] .power_up = "low";

dffeas \out_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[46]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_46),
	.prn(vcc));
defparam \out_data_buffer[46] .is_wysiwyg = "true";
defparam \out_data_buffer[46] .power_up = "low";

dffeas \out_data_buffer[47] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[47]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_47),
	.prn(vcc));
defparam \out_data_buffer[47] .is_wysiwyg = "true";
defparam \out_data_buffer[47] .power_up = "low";

dffeas \out_data_buffer[32] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[32]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_32),
	.prn(vcc));
defparam \out_data_buffer[32] .is_wysiwyg = "true";
defparam \out_data_buffer[32] .power_up = "low";

dffeas \out_data_buffer[33] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[33]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_33),
	.prn(vcc));
defparam \out_data_buffer[33] .is_wysiwyg = "true";
defparam \out_data_buffer[33] .power_up = "low";

dffeas \out_data_buffer[34] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[34]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_34),
	.prn(vcc));
defparam \out_data_buffer[34] .is_wysiwyg = "true";
defparam \out_data_buffer[34] .power_up = "low";

dffeas \out_data_buffer[35] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[35]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_35),
	.prn(vcc));
defparam \out_data_buffer[35] .is_wysiwyg = "true";
defparam \out_data_buffer[35] .power_up = "low";

cycloneive_lcell_comb \take_in_data~2 (
	.dataa(Equal1),
	.datab(always1),
	.datac(Equal2),
	.datad(\in_ready~0_combout ),
	.cin(gnd),
	.combout(take_in_data),
	.cout());
defparam \take_in_data~2 .lut_mask = 16'hBFFF;
defparam \take_in_data~2 .sum_lutc_input = "datac";

dffeas \out_data_buffer[107] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[107]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_107),
	.prn(vcc));
defparam \out_data_buffer[107] .is_wysiwyg = "true";
defparam \out_data_buffer[107] .power_up = "low";

dffeas \out_data_buffer[86] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[86]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_86),
	.prn(vcc));
defparam \out_data_buffer[86] .is_wysiwyg = "true";
defparam \out_data_buffer[86] .power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(\in_to_out_synchronizer|dreg[0]~q ),
	.datab(\out_data_toggle_flopped~q ),
	.datac(last_cycle),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_toggle_flopped~q ),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb \take_in_data~3 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(take_in_data),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~3_combout ),
	.cout());
defparam \take_in_data~3 .lut_mask = 16'hF7F7;
defparam \take_in_data~3 .sum_lutc_input = "datac";

dffeas \in_data_buffer[68] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[68]~q ),
	.prn(vcc));
defparam \in_data_buffer[68] .is_wysiwyg = "true";
defparam \in_data_buffer[68] .power_up = "low";

dffeas \in_data_buffer[48] (
	.clk(clk_clk),
	.d(in_data[48]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[48]~q ),
	.prn(vcc));
defparam \in_data_buffer[48] .is_wysiwyg = "true";
defparam \in_data_buffer[48] .power_up = "low";

dffeas \in_data_buffer[62] (
	.clk(clk_clk),
	.d(in_data[62]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[62]~q ),
	.prn(vcc));
defparam \in_data_buffer[62] .is_wysiwyg = "true";
defparam \in_data_buffer[62] .power_up = "low";

dffeas \in_data_buffer[49] (
	.clk(clk_clk),
	.d(in_data[49]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[49]~q ),
	.prn(vcc));
defparam \in_data_buffer[49] .is_wysiwyg = "true";
defparam \in_data_buffer[49] .power_up = "low";

dffeas \in_data_buffer[51] (
	.clk(clk_clk),
	.d(in_data[51]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[51]~q ),
	.prn(vcc));
defparam \in_data_buffer[51] .is_wysiwyg = "true";
defparam \in_data_buffer[51] .power_up = "low";

dffeas \in_data_buffer[50] (
	.clk(clk_clk),
	.d(in_data[50]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[50]~q ),
	.prn(vcc));
defparam \in_data_buffer[50] .is_wysiwyg = "true";
defparam \in_data_buffer[50] .power_up = "low";

dffeas \in_data_buffer[53] (
	.clk(clk_clk),
	.d(in_data[53]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[53]~q ),
	.prn(vcc));
defparam \in_data_buffer[53] .is_wysiwyg = "true";
defparam \in_data_buffer[53] .power_up = "low";

dffeas \in_data_buffer[52] (
	.clk(clk_clk),
	.d(in_data[52]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[52]~q ),
	.prn(vcc));
defparam \in_data_buffer[52] .is_wysiwyg = "true";
defparam \in_data_buffer[52] .power_up = "low";

dffeas \in_data_buffer[55] (
	.clk(clk_clk),
	.d(in_data[55]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[55]~q ),
	.prn(vcc));
defparam \in_data_buffer[55] .is_wysiwyg = "true";
defparam \in_data_buffer[55] .power_up = "low";

dffeas \in_data_buffer[54] (
	.clk(clk_clk),
	.d(in_data[54]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[54]~q ),
	.prn(vcc));
defparam \in_data_buffer[54] .is_wysiwyg = "true";
defparam \in_data_buffer[54] .power_up = "low";

dffeas \in_data_buffer[57] (
	.clk(clk_clk),
	.d(in_data[57]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[57]~q ),
	.prn(vcc));
defparam \in_data_buffer[57] .is_wysiwyg = "true";
defparam \in_data_buffer[57] .power_up = "low";

dffeas \in_data_buffer[56] (
	.clk(clk_clk),
	.d(in_data[56]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[56]~q ),
	.prn(vcc));
defparam \in_data_buffer[56] .is_wysiwyg = "true";
defparam \in_data_buffer[56] .power_up = "low";

dffeas \in_data_buffer[59] (
	.clk(clk_clk),
	.d(in_data[59]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[59]~q ),
	.prn(vcc));
defparam \in_data_buffer[59] .is_wysiwyg = "true";
defparam \in_data_buffer[59] .power_up = "low";

dffeas \in_data_buffer[58] (
	.clk(clk_clk),
	.d(in_data[58]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[58]~q ),
	.prn(vcc));
defparam \in_data_buffer[58] .is_wysiwyg = "true";
defparam \in_data_buffer[58] .power_up = "low";

dffeas \in_data_buffer[61] (
	.clk(clk_clk),
	.d(in_data[61]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[61]~q ),
	.prn(vcc));
defparam \in_data_buffer[61] .is_wysiwyg = "true";
defparam \in_data_buffer[61] .power_up = "low";

dffeas \in_data_buffer[60] (
	.clk(clk_clk),
	.d(in_data[60]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[60]~q ),
	.prn(vcc));
defparam \in_data_buffer[60] .is_wysiwyg = "true";
defparam \in_data_buffer[60] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(clk_clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(clk_clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[40] (
	.clk(clk_clk),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[40]~q ),
	.prn(vcc));
defparam \in_data_buffer[40] .is_wysiwyg = "true";
defparam \in_data_buffer[40] .power_up = "low";

dffeas \in_data_buffer[41] (
	.clk(clk_clk),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[41]~q ),
	.prn(vcc));
defparam \in_data_buffer[41] .is_wysiwyg = "true";
defparam \in_data_buffer[41] .power_up = "low";

dffeas \in_data_buffer[42] (
	.clk(clk_clk),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[42]~q ),
	.prn(vcc));
defparam \in_data_buffer[42] .is_wysiwyg = "true";
defparam \in_data_buffer[42] .power_up = "low";

dffeas \in_data_buffer[43] (
	.clk(clk_clk),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[43]~q ),
	.prn(vcc));
defparam \in_data_buffer[43] .is_wysiwyg = "true";
defparam \in_data_buffer[43] .power_up = "low";

dffeas \in_data_buffer[44] (
	.clk(clk_clk),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[44]~q ),
	.prn(vcc));
defparam \in_data_buffer[44] .is_wysiwyg = "true";
defparam \in_data_buffer[44] .power_up = "low";

dffeas \in_data_buffer[45] (
	.clk(clk_clk),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[45]~q ),
	.prn(vcc));
defparam \in_data_buffer[45] .is_wysiwyg = "true";
defparam \in_data_buffer[45] .power_up = "low";

dffeas \in_data_buffer[46] (
	.clk(clk_clk),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[46]~q ),
	.prn(vcc));
defparam \in_data_buffer[46] .is_wysiwyg = "true";
defparam \in_data_buffer[46] .power_up = "low";

dffeas \in_data_buffer[47] (
	.clk(clk_clk),
	.d(in_data[47]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[47]~q ),
	.prn(vcc));
defparam \in_data_buffer[47] .is_wysiwyg = "true";
defparam \in_data_buffer[47] .power_up = "low";

dffeas \in_data_buffer[32] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[32]~q ),
	.prn(vcc));
defparam \in_data_buffer[32] .is_wysiwyg = "true";
defparam \in_data_buffer[32] .power_up = "low";

dffeas \in_data_buffer[33] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[33]~q ),
	.prn(vcc));
defparam \in_data_buffer[33] .is_wysiwyg = "true";
defparam \in_data_buffer[33] .power_up = "low";

dffeas \in_data_buffer[34] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[34]~q ),
	.prn(vcc));
defparam \in_data_buffer[34] .is_wysiwyg = "true";
defparam \in_data_buffer[34] .power_up = "low";

dffeas \in_data_buffer[35] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[35]~q ),
	.prn(vcc));
defparam \in_data_buffer[35] .is_wysiwyg = "true";
defparam \in_data_buffer[35] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(\in_data_toggle~q ),
	.datad(take_in_data),
	.cin(gnd),
	.combout(\in_data_toggle~2_combout ),
	.cout());
defparam \in_data_toggle~2 .lut_mask = 16'h6996;
defparam \in_data_toggle~2 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~2_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \in_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\in_ready~0_combout ),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h0FF0;
defparam \in_ready~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[107] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[107]~q ),
	.prn(vcc));
defparam \in_data_buffer[107] .is_wysiwyg = "true";
defparam \in_data_buffer[107] .power_up = "low";

dffeas \in_data_buffer[86] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~3_combout ),
	.q(\in_data_buffer[86]~q ),
	.prn(vcc));
defparam \in_data_buffer[86] .is_wysiwyg = "true";
defparam \in_data_buffer[86] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_6 (
	clk,
	reset_n,
	dreg_0,
	din)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	dreg_0;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_7 (
	reset_n,
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_avalon_st_handshake_clock_crosser_2 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_buffer_67,
	mem_used_0,
	mem_107_0,
	out_valid1,
	in_data_toggle,
	dreg_01,
	always0,
	out_data_buffer_0,
	mem_67_0,
	take_in_data,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_18,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_24,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_22,
	out_payload_23,
	out_payload_24,
	out_payload_25,
	out_payload_26,
	out_payload_11,
	out_payload_13,
	out_payload_16,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_10,
	out_payload_9,
	out_payload_8,
	out_payload_7,
	out_payload_6,
	out_payload_20,
	out_payload_18,
	out_payload_19,
	out_payload_17,
	out_payload_21,
	out_data_buffer_31,
	out_payload_27,
	out_data_buffer_30,
	out_data_buffer_29,
	out_payload_28,
	out_payload_31,
	out_payload_30,
	out_payload_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
output 	out_data_buffer_67;
input 	mem_used_0;
input 	mem_107_0;
input 	out_valid1;
output 	in_data_toggle;
output 	dreg_01;
input 	always0;
output 	out_data_buffer_0;
input 	mem_67_0;
output 	take_in_data;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_18;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_24;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
input 	out_payload_0;
input 	out_payload_1;
input 	out_payload_2;
input 	out_payload_3;
input 	out_payload_4;
input 	out_payload_22;
input 	out_payload_23;
input 	out_payload_24;
input 	out_payload_25;
input 	out_payload_26;
input 	out_payload_11;
input 	out_payload_13;
input 	out_payload_16;
input 	out_payload_12;
input 	out_payload_5;
input 	out_payload_14;
input 	out_payload_15;
input 	out_payload_10;
input 	out_payload_9;
input 	out_payload_8;
input 	out_payload_7;
input 	out_payload_6;
input 	out_payload_20;
input 	out_payload_18;
input 	out_payload_19;
input 	out_payload_17;
input 	out_payload_21;
output 	out_data_buffer_31;
input 	out_payload_27;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
input 	out_payload_28;
input 	out_payload_31;
input 	out_payload_30;
input 	out_payload_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_avalon_st_clock_crosser_1 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.mem_used_0(mem_used_0),
	.mem_107_0(mem_107_0),
	.out_valid2(out_valid1),
	.in_data_toggle1(in_data_toggle),
	.dreg_01(dreg_01),
	.always0(always0),
	.out_data_buffer_0(out_data_buffer_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,mem_67_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_payload_31,out_payload_30,out_payload_29,out_payload_28,out_payload_27,out_payload_26,out_payload_25,out_payload_24,out_payload_23,out_payload_22,out_payload_21,out_payload_20,out_payload_19,out_payload_18,out_payload_17,out_payload_16,out_payload_15,
out_payload_14,out_payload_13,out_payload_12,out_payload_11,out_payload_10,out_payload_9,out_payload_8,out_payload_7,out_payload_6,out_payload_5,out_payload_4,out_payload_3,out_payload_2,out_payload_1,out_payload_0}),
	.take_in_data(take_in_data),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.clk_clk(clk_clk));

endmodule

module usb_system_altera_avalon_st_clock_crosser_1 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	out_data_buffer_67,
	mem_used_0,
	mem_107_0,
	out_valid2,
	in_data_toggle1,
	dreg_01,
	always0,
	out_data_buffer_0,
	in_data,
	take_in_data,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_18,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_24,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
output 	out_data_buffer_67;
input 	mem_used_0;
input 	mem_107_0;
input 	out_valid2;
output 	in_data_toggle1;
output 	dreg_01;
input 	always0;
output 	out_data_buffer_0;
input 	[118:0] in_data;
output 	take_in_data;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_18;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_24;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \take_in_data~1_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;


usb_system_altera_std_synchronizer_9 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(dreg_01));

usb_system_altera_std_synchronizer_8 in_to_out_synchronizer(
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(in_data_toggle1),
	.clk(clk_clk));

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_clk),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(out_valid2),
	.datab(mem_used_0),
	.datac(mem_107_0),
	.datad(gnd),
	.cin(gnd),
	.combout(take_in_data),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hFEFE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_clk),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_clk),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(clk_clk),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_clk),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_clk),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_clk),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_clk),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_clk),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_clk),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_clk),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_clk),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_clk),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_clk),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_clk),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_clk),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_clk),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_clk),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_clk),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_clk),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_clk),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_clk),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_clk),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_clk),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

cycloneive_lcell_comb \take_in_data~1 (
	.dataa(take_in_data),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(always0),
	.cin(gnd),
	.combout(\take_in_data~1_combout ),
	.cout());
defparam \take_in_data~1 .lut_mask = 16'hBEFF;
defparam \take_in_data~1 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(wire_pll7_clk_0),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(always0),
	.datac(take_in_data),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_8 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_9 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_avalon_st_handshake_clock_crosser_3 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_buffer_67,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	in_data_toggle,
	dreg_01,
	always0,
	out_data_buffer_22,
	out_data_buffer_23,
	out_data_buffer_24,
	out_data_buffer_25,
	out_data_buffer_26,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_20,
	out_data_buffer_18,
	out_data_buffer_19,
	out_data_buffer_17,
	out_data_buffer_21,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	mem_67_0,
	take_in_data,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_22,
	out_payload_23,
	out_payload_24,
	out_payload_25,
	out_payload_26,
	out_payload_11,
	out_payload_13,
	out_payload_16,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_10,
	out_payload_9,
	out_payload_8,
	out_payload_7,
	out_payload_6,
	out_payload_20,
	out_payload_18,
	out_payload_19,
	out_payload_17,
	out_payload_21,
	out_payload_27,
	out_payload_28,
	out_payload_31,
	out_payload_30,
	out_payload_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
output 	out_data_buffer_67;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	in_data_toggle;
output 	dreg_01;
input 	always0;
output 	out_data_buffer_22;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_20;
output 	out_data_buffer_18;
output 	out_data_buffer_19;
output 	out_data_buffer_17;
output 	out_data_buffer_21;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
input 	mem_67_0;
input 	take_in_data;
input 	out_payload_0;
input 	out_payload_1;
input 	out_payload_2;
input 	out_payload_3;
input 	out_payload_4;
input 	out_payload_22;
input 	out_payload_23;
input 	out_payload_24;
input 	out_payload_25;
input 	out_payload_26;
input 	out_payload_11;
input 	out_payload_13;
input 	out_payload_16;
input 	out_payload_12;
input 	out_payload_5;
input 	out_payload_14;
input 	out_payload_15;
input 	out_payload_10;
input 	out_payload_9;
input 	out_payload_8;
input 	out_payload_7;
input 	out_payload_6;
input 	out_payload_20;
input 	out_payload_18;
input 	out_payload_19;
input 	out_payload_17;
input 	out_payload_21;
input 	out_payload_27;
input 	out_payload_28;
input 	out_payload_31;
input 	out_payload_30;
input 	out_payload_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_avalon_st_clock_crosser_2 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.in_data_toggle1(in_data_toggle),
	.dreg_01(dreg_01),
	.always0(always0),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,mem_67_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_payload_31,out_payload_30,out_payload_29,out_payload_28,out_payload_27,out_payload_26,out_payload_25,out_payload_24,out_payload_23,out_payload_22,out_payload_21,out_payload_20,out_payload_19,out_payload_18,out_payload_17,out_payload_16,out_payload_15,
out_payload_14,out_payload_13,out_payload_12,out_payload_11,out_payload_10,out_payload_9,out_payload_8,out_payload_7,out_payload_6,out_payload_5,out_payload_4,out_payload_3,out_payload_2,out_payload_1,out_payload_0}),
	.take_in_data(take_in_data),
	.clk_clk(clk_clk));

endmodule

module usb_system_altera_avalon_st_clock_crosser_2 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	out_data_buffer_67,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	in_data_toggle1,
	dreg_01,
	always0,
	out_data_buffer_22,
	out_data_buffer_23,
	out_data_buffer_24,
	out_data_buffer_25,
	out_data_buffer_26,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_20,
	out_data_buffer_18,
	out_data_buffer_19,
	out_data_buffer_17,
	out_data_buffer_21,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	in_data,
	take_in_data,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
output 	out_data_buffer_67;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	in_data_toggle1;
output 	dreg_01;
input 	always0;
output 	out_data_buffer_22;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_20;
output 	out_data_buffer_18;
output 	out_data_buffer_19;
output 	out_data_buffer_17;
output 	out_data_buffer_21;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
input 	[118:0] in_data;
input 	take_in_data;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \take_in_data~0_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;


usb_system_altera_std_synchronizer_11 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(dreg_01));

usb_system_altera_std_synchronizer_10 in_to_out_synchronizer(
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(in_data_toggle1),
	.clk(clk_clk));

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_clk),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_clk),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_clk),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_clk),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_clk),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_clk),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(clk_clk),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_clk),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_clk),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_clk),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_clk),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_clk),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_clk),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_clk),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_clk),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_clk),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_clk),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_clk),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_clk),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_clk),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_clk),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_clk),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_clk),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_clk),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(always0),
	.datab(take_in_data),
	.datac(in_data_toggle1),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\take_in_data~0_combout ),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hEFFE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(wire_pll7_clk_0),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(always0),
	.datac(take_in_data),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_10 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_11 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_avalon_st_clock_crosser_3 (
	wire_pll7_clk_0,
	in_data,
	in_reset,
	out_reset,
	sink_ready,
	in_data_toggle1,
	dreg_0,
	s0_cmd_valid,
	last_cycle,
	saved_grant_0,
	out_data_toggle_flopped1,
	dreg_01,
	out_valid1,
	out_data_buffer_67,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	sink_ready1,
	out_data_buffer_107,
	out_data_buffer_66,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_18,
	out_data_buffer_19,
	out_data_buffer_20,
	out_data_buffer_21,
	out_data_buffer_22,
	out_data_buffer_23,
	out_data_buffer_24,
	out_data_buffer_25,
	out_data_buffer_26,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_29,
	out_data_buffer_30,
	out_data_buffer_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	[118:0] in_data;
input 	in_reset;
input 	out_reset;
input 	sink_ready;
output 	in_data_toggle1;
output 	dreg_0;
input 	s0_cmd_valid;
input 	last_cycle;
input 	saved_grant_0;
output 	out_data_toggle_flopped1;
output 	dreg_01;
output 	out_valid1;
output 	out_data_buffer_67;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
input 	sink_ready1;
output 	out_data_buffer_107;
output 	out_data_buffer_66;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_18;
output 	out_data_buffer_19;
output 	out_data_buffer_20;
output 	out_data_buffer_21;
output 	out_data_buffer_22;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_29;
output 	out_data_buffer_30;
output 	out_data_buffer_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_data_toggle~0_combout ;
wire \out_data_toggle_flopped~0_combout ;
wire \take_in_data~combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_buffer[68]~q ;
wire \in_data_buffer[48]~q ;
wire \in_data_buffer[62]~q ;
wire \in_data_buffer[49]~q ;
wire \in_data_buffer[51]~q ;
wire \in_data_buffer[50]~q ;
wire \in_data_buffer[53]~q ;
wire \in_data_buffer[52]~q ;
wire \in_data_buffer[55]~q ;
wire \in_data_buffer[54]~q ;
wire \in_data_buffer[57]~q ;
wire \in_data_buffer[56]~q ;
wire \in_data_buffer[59]~q ;
wire \in_data_buffer[58]~q ;
wire \in_data_buffer[61]~q ;
wire \in_data_buffer[60]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[40]~q ;
wire \in_data_buffer[41]~q ;
wire \in_data_buffer[42]~q ;
wire \in_data_buffer[43]~q ;
wire \in_data_buffer[44]~q ;
wire \in_data_buffer[45]~q ;
wire \in_data_buffer[46]~q ;
wire \in_data_buffer[47]~q ;
wire \in_data_buffer[32]~q ;
wire \in_data_buffer[33]~q ;
wire \in_data_buffer[34]~q ;
wire \in_data_buffer[35]~q ;
wire \in_data_buffer[107]~q ;
wire \in_data_buffer[66]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[31]~q ;


usb_system_altera_std_synchronizer_13 out_to_in_synchronizer(
	.reset_n(in_reset),
	.dreg_0(dreg_0),
	.din(out_data_toggle_flopped1),
	.clk(clk_clk));

usb_system_altera_std_synchronizer_12 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.din(in_data_toggle1),
	.dreg_0(dreg_01));

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_01),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas \out_data_buffer[68] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[68]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_68),
	.prn(vcc));
defparam \out_data_buffer[68] .is_wysiwyg = "true";
defparam \out_data_buffer[68] .power_up = "low";

dffeas \out_data_buffer[48] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[48]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_48),
	.prn(vcc));
defparam \out_data_buffer[48] .is_wysiwyg = "true";
defparam \out_data_buffer[48] .power_up = "low";

dffeas \out_data_buffer[62] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[62]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_62),
	.prn(vcc));
defparam \out_data_buffer[62] .is_wysiwyg = "true";
defparam \out_data_buffer[62] .power_up = "low";

dffeas \out_data_buffer[49] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[49]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_49),
	.prn(vcc));
defparam \out_data_buffer[49] .is_wysiwyg = "true";
defparam \out_data_buffer[49] .power_up = "low";

dffeas \out_data_buffer[51] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[51]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_51),
	.prn(vcc));
defparam \out_data_buffer[51] .is_wysiwyg = "true";
defparam \out_data_buffer[51] .power_up = "low";

dffeas \out_data_buffer[50] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[50]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_50),
	.prn(vcc));
defparam \out_data_buffer[50] .is_wysiwyg = "true";
defparam \out_data_buffer[50] .power_up = "low";

dffeas \out_data_buffer[53] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[53]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_53),
	.prn(vcc));
defparam \out_data_buffer[53] .is_wysiwyg = "true";
defparam \out_data_buffer[53] .power_up = "low";

dffeas \out_data_buffer[52] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[52]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_52),
	.prn(vcc));
defparam \out_data_buffer[52] .is_wysiwyg = "true";
defparam \out_data_buffer[52] .power_up = "low";

dffeas \out_data_buffer[55] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[55]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_55),
	.prn(vcc));
defparam \out_data_buffer[55] .is_wysiwyg = "true";
defparam \out_data_buffer[55] .power_up = "low";

dffeas \out_data_buffer[54] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[54]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_54),
	.prn(vcc));
defparam \out_data_buffer[54] .is_wysiwyg = "true";
defparam \out_data_buffer[54] .power_up = "low";

dffeas \out_data_buffer[57] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[57]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_57),
	.prn(vcc));
defparam \out_data_buffer[57] .is_wysiwyg = "true";
defparam \out_data_buffer[57] .power_up = "low";

dffeas \out_data_buffer[56] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[56]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_56),
	.prn(vcc));
defparam \out_data_buffer[56] .is_wysiwyg = "true";
defparam \out_data_buffer[56] .power_up = "low";

dffeas \out_data_buffer[59] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[59]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_59),
	.prn(vcc));
defparam \out_data_buffer[59] .is_wysiwyg = "true";
defparam \out_data_buffer[59] .power_up = "low";

dffeas \out_data_buffer[58] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[58]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_58),
	.prn(vcc));
defparam \out_data_buffer[58] .is_wysiwyg = "true";
defparam \out_data_buffer[58] .power_up = "low";

dffeas \out_data_buffer[61] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[61]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_61),
	.prn(vcc));
defparam \out_data_buffer[61] .is_wysiwyg = "true";
defparam \out_data_buffer[61] .power_up = "low";

dffeas \out_data_buffer[60] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[60]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_60),
	.prn(vcc));
defparam \out_data_buffer[60] .is_wysiwyg = "true";
defparam \out_data_buffer[60] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas \out_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[40]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_40),
	.prn(vcc));
defparam \out_data_buffer[40] .is_wysiwyg = "true";
defparam \out_data_buffer[40] .power_up = "low";

dffeas \out_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[41]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_41),
	.prn(vcc));
defparam \out_data_buffer[41] .is_wysiwyg = "true";
defparam \out_data_buffer[41] .power_up = "low";

dffeas \out_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[42]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_42),
	.prn(vcc));
defparam \out_data_buffer[42] .is_wysiwyg = "true";
defparam \out_data_buffer[42] .power_up = "low";

dffeas \out_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[43]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_43),
	.prn(vcc));
defparam \out_data_buffer[43] .is_wysiwyg = "true";
defparam \out_data_buffer[43] .power_up = "low";

dffeas \out_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[44]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_44),
	.prn(vcc));
defparam \out_data_buffer[44] .is_wysiwyg = "true";
defparam \out_data_buffer[44] .power_up = "low";

dffeas \out_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[45]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_45),
	.prn(vcc));
defparam \out_data_buffer[45] .is_wysiwyg = "true";
defparam \out_data_buffer[45] .power_up = "low";

dffeas \out_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[46]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_46),
	.prn(vcc));
defparam \out_data_buffer[46] .is_wysiwyg = "true";
defparam \out_data_buffer[46] .power_up = "low";

dffeas \out_data_buffer[47] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[47]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_47),
	.prn(vcc));
defparam \out_data_buffer[47] .is_wysiwyg = "true";
defparam \out_data_buffer[47] .power_up = "low";

dffeas \out_data_buffer[32] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[32]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_32),
	.prn(vcc));
defparam \out_data_buffer[32] .is_wysiwyg = "true";
defparam \out_data_buffer[32] .power_up = "low";

dffeas \out_data_buffer[33] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[33]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_33),
	.prn(vcc));
defparam \out_data_buffer[33] .is_wysiwyg = "true";
defparam \out_data_buffer[33] .power_up = "low";

dffeas \out_data_buffer[34] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[34]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_34),
	.prn(vcc));
defparam \out_data_buffer[34] .is_wysiwyg = "true";
defparam \out_data_buffer[34] .power_up = "low";

dffeas \out_data_buffer[35] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[35]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_35),
	.prn(vcc));
defparam \out_data_buffer[35] .is_wysiwyg = "true";
defparam \out_data_buffer[35] .power_up = "low";

dffeas \out_data_buffer[107] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[107]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_107),
	.prn(vcc));
defparam \out_data_buffer[107] .is_wysiwyg = "true";
defparam \out_data_buffer[107] .power_up = "low";

dffeas \out_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(sink_ready),
	.datac(sink_ready1),
	.datad(s0_cmd_valid),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'h6996;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(dreg_01),
	.datab(out_data_toggle_flopped1),
	.datac(last_cycle),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb take_in_data(
	.dataa(sink_ready),
	.datab(sink_ready1),
	.datac(s0_cmd_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hFEFE;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(clk_clk),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

dffeas \in_data_buffer[68] (
	.clk(clk_clk),
	.d(in_data[68]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[68]~q ),
	.prn(vcc));
defparam \in_data_buffer[68] .is_wysiwyg = "true";
defparam \in_data_buffer[68] .power_up = "low";

dffeas \in_data_buffer[48] (
	.clk(clk_clk),
	.d(in_data[48]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[48]~q ),
	.prn(vcc));
defparam \in_data_buffer[48] .is_wysiwyg = "true";
defparam \in_data_buffer[48] .power_up = "low";

dffeas \in_data_buffer[62] (
	.clk(clk_clk),
	.d(in_data[62]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[62]~q ),
	.prn(vcc));
defparam \in_data_buffer[62] .is_wysiwyg = "true";
defparam \in_data_buffer[62] .power_up = "low";

dffeas \in_data_buffer[49] (
	.clk(clk_clk),
	.d(in_data[49]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[49]~q ),
	.prn(vcc));
defparam \in_data_buffer[49] .is_wysiwyg = "true";
defparam \in_data_buffer[49] .power_up = "low";

dffeas \in_data_buffer[51] (
	.clk(clk_clk),
	.d(in_data[51]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[51]~q ),
	.prn(vcc));
defparam \in_data_buffer[51] .is_wysiwyg = "true";
defparam \in_data_buffer[51] .power_up = "low";

dffeas \in_data_buffer[50] (
	.clk(clk_clk),
	.d(in_data[50]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[50]~q ),
	.prn(vcc));
defparam \in_data_buffer[50] .is_wysiwyg = "true";
defparam \in_data_buffer[50] .power_up = "low";

dffeas \in_data_buffer[53] (
	.clk(clk_clk),
	.d(in_data[53]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[53]~q ),
	.prn(vcc));
defparam \in_data_buffer[53] .is_wysiwyg = "true";
defparam \in_data_buffer[53] .power_up = "low";

dffeas \in_data_buffer[52] (
	.clk(clk_clk),
	.d(in_data[52]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[52]~q ),
	.prn(vcc));
defparam \in_data_buffer[52] .is_wysiwyg = "true";
defparam \in_data_buffer[52] .power_up = "low";

dffeas \in_data_buffer[55] (
	.clk(clk_clk),
	.d(in_data[55]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[55]~q ),
	.prn(vcc));
defparam \in_data_buffer[55] .is_wysiwyg = "true";
defparam \in_data_buffer[55] .power_up = "low";

dffeas \in_data_buffer[54] (
	.clk(clk_clk),
	.d(in_data[54]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[54]~q ),
	.prn(vcc));
defparam \in_data_buffer[54] .is_wysiwyg = "true";
defparam \in_data_buffer[54] .power_up = "low";

dffeas \in_data_buffer[57] (
	.clk(clk_clk),
	.d(in_data[57]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[57]~q ),
	.prn(vcc));
defparam \in_data_buffer[57] .is_wysiwyg = "true";
defparam \in_data_buffer[57] .power_up = "low";

dffeas \in_data_buffer[56] (
	.clk(clk_clk),
	.d(in_data[56]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[56]~q ),
	.prn(vcc));
defparam \in_data_buffer[56] .is_wysiwyg = "true";
defparam \in_data_buffer[56] .power_up = "low";

dffeas \in_data_buffer[59] (
	.clk(clk_clk),
	.d(in_data[59]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[59]~q ),
	.prn(vcc));
defparam \in_data_buffer[59] .is_wysiwyg = "true";
defparam \in_data_buffer[59] .power_up = "low";

dffeas \in_data_buffer[58] (
	.clk(clk_clk),
	.d(in_data[58]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[58]~q ),
	.prn(vcc));
defparam \in_data_buffer[58] .is_wysiwyg = "true";
defparam \in_data_buffer[58] .power_up = "low";

dffeas \in_data_buffer[61] (
	.clk(clk_clk),
	.d(in_data[61]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[61]~q ),
	.prn(vcc));
defparam \in_data_buffer[61] .is_wysiwyg = "true";
defparam \in_data_buffer[61] .power_up = "low";

dffeas \in_data_buffer[60] (
	.clk(clk_clk),
	.d(in_data[60]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[60]~q ),
	.prn(vcc));
defparam \in_data_buffer[60] .is_wysiwyg = "true";
defparam \in_data_buffer[60] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(clk_clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(clk_clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[40] (
	.clk(clk_clk),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[40]~q ),
	.prn(vcc));
defparam \in_data_buffer[40] .is_wysiwyg = "true";
defparam \in_data_buffer[40] .power_up = "low";

dffeas \in_data_buffer[41] (
	.clk(clk_clk),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[41]~q ),
	.prn(vcc));
defparam \in_data_buffer[41] .is_wysiwyg = "true";
defparam \in_data_buffer[41] .power_up = "low";

dffeas \in_data_buffer[42] (
	.clk(clk_clk),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[42]~q ),
	.prn(vcc));
defparam \in_data_buffer[42] .is_wysiwyg = "true";
defparam \in_data_buffer[42] .power_up = "low";

dffeas \in_data_buffer[43] (
	.clk(clk_clk),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[43]~q ),
	.prn(vcc));
defparam \in_data_buffer[43] .is_wysiwyg = "true";
defparam \in_data_buffer[43] .power_up = "low";

dffeas \in_data_buffer[44] (
	.clk(clk_clk),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[44]~q ),
	.prn(vcc));
defparam \in_data_buffer[44] .is_wysiwyg = "true";
defparam \in_data_buffer[44] .power_up = "low";

dffeas \in_data_buffer[45] (
	.clk(clk_clk),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[45]~q ),
	.prn(vcc));
defparam \in_data_buffer[45] .is_wysiwyg = "true";
defparam \in_data_buffer[45] .power_up = "low";

dffeas \in_data_buffer[46] (
	.clk(clk_clk),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[46]~q ),
	.prn(vcc));
defparam \in_data_buffer[46] .is_wysiwyg = "true";
defparam \in_data_buffer[46] .power_up = "low";

dffeas \in_data_buffer[47] (
	.clk(clk_clk),
	.d(in_data[47]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[47]~q ),
	.prn(vcc));
defparam \in_data_buffer[47] .is_wysiwyg = "true";
defparam \in_data_buffer[47] .power_up = "low";

dffeas \in_data_buffer[32] (
	.clk(clk_clk),
	.d(in_data[32]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[32]~q ),
	.prn(vcc));
defparam \in_data_buffer[32] .is_wysiwyg = "true";
defparam \in_data_buffer[32] .power_up = "low";

dffeas \in_data_buffer[33] (
	.clk(clk_clk),
	.d(in_data[33]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[33]~q ),
	.prn(vcc));
defparam \in_data_buffer[33] .is_wysiwyg = "true";
defparam \in_data_buffer[33] .power_up = "low";

dffeas \in_data_buffer[34] (
	.clk(clk_clk),
	.d(in_data[34]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[34]~q ),
	.prn(vcc));
defparam \in_data_buffer[34] .is_wysiwyg = "true";
defparam \in_data_buffer[34] .power_up = "low";

dffeas \in_data_buffer[35] (
	.clk(clk_clk),
	.d(in_data[35]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[35]~q ),
	.prn(vcc));
defparam \in_data_buffer[35] .is_wysiwyg = "true";
defparam \in_data_buffer[35] .power_up = "low";

dffeas \in_data_buffer[107] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[107]~q ),
	.prn(vcc));
defparam \in_data_buffer[107] .is_wysiwyg = "true";
defparam \in_data_buffer[107] .power_up = "low";

dffeas \in_data_buffer[66] (
	.clk(clk_clk),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(clk_clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(clk_clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(clk_clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(clk_clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(clk_clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(clk_clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(clk_clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(clk_clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(clk_clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(clk_clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(clk_clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(clk_clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(clk_clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(clk_clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(clk_clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(clk_clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(clk_clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(clk_clk),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(clk_clk),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(clk_clk),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(clk_clk),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(clk_clk),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(clk_clk),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(clk_clk),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(clk_clk),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(clk_clk),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_12 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_std_synchronizer_13 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module usb_system_altera_merlin_master_agent_1 (
	mem_67_0,
	mem_67_01,
	mem_67_02,
	src1_valid,
	src_payload,
	out_valid,
	src_payload1,
	WideOr1,
	av_readdatavalid,
	out_data_buffer_67,
	av_readdatavalid1,
	av_readdatavalid2)/* synthesis synthesis_greybox=1 */;
input 	mem_67_0;
input 	mem_67_01;
input 	mem_67_02;
input 	src1_valid;
input 	src_payload;
input 	out_valid;
input 	src_payload1;
input 	WideOr1;
output 	av_readdatavalid;
input 	out_data_buffer_67;
output 	av_readdatavalid1;
output 	av_readdatavalid2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \av_readdatavalid~0 (
	.dataa(mem_67_0),
	.datab(src_payload1),
	.datac(mem_67_02),
	.datad(src_payload),
	.cin(gnd),
	.combout(av_readdatavalid),
	.cout());
defparam \av_readdatavalid~0 .lut_mask = 16'h7FFF;
defparam \av_readdatavalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdatavalid~1 (
	.dataa(mem_67_01),
	.datab(src1_valid),
	.datac(out_valid),
	.datad(out_data_buffer_67),
	.cin(gnd),
	.combout(av_readdatavalid1),
	.cout());
defparam \av_readdatavalid~1 .lut_mask = 16'h7FFF;
defparam \av_readdatavalid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdatavalid~2 (
	.dataa(WideOr1),
	.datab(av_readdatavalid),
	.datac(av_readdatavalid1),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdatavalid2),
	.cout());
defparam \av_readdatavalid~2 .lut_mask = 16'hFEFE;
defparam \av_readdatavalid~2 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_master_translator (
	reset,
	d_write,
	write_accepted1,
	sink_in_reset,
	d_read,
	read_accepted1,
	av_ld_getting_data,
	uav_write,
	uav_read,
	WideOr0,
	av_waitrequest,
	s0_cmd_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
output 	write_accepted1;
input 	sink_in_reset;
input 	d_read;
output 	read_accepted1;
input 	av_ld_getting_data;
output 	uav_write;
output 	uav_read;
input 	WideOr0;
output 	av_waitrequest;
input 	s0_cmd_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write_accepted~0_combout ;
wire \write_accepted~1_combout ;
wire \read_accepted~0_combout ;
wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;
wire \av_waitrequest~0_combout ;


dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb \uav_write~0 (
	.dataa(d_write),
	.datab(gnd),
	.datac(gnd),
	.datad(write_accepted1),
	.cin(gnd),
	.combout(uav_write),
	.cout());
defparam \uav_write~0 .lut_mask = 16'hAAFF;
defparam \uav_write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \uav_read~0 (
	.dataa(d_read),
	.datab(gnd),
	.datac(gnd),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read),
	.cout());
defparam \uav_read~0 .lut_mask = 16'hAAFF;
defparam \uav_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~1 (
	.dataa(d_read),
	.datab(d_write),
	.datac(av_ld_getting_data),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(av_waitrequest),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'h27FF;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_accepted~0 (
	.dataa(sink_in_reset),
	.datab(WideOr0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_accepted~0_combout ),
	.cout());
defparam \write_accepted~0 .lut_mask = 16'hEEEE;
defparam \write_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_accepted~1 (
	.dataa(av_waitrequest),
	.datab(write_accepted1),
	.datac(d_write),
	.datad(\write_accepted~0_combout ),
	.cin(gnd),
	.combout(\write_accepted~1_combout ),
	.cout());
defparam \write_accepted~1 .lut_mask = 16'hFFFE;
defparam \write_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(read_accepted1),
	.datab(d_read),
	.datac(\write_accepted~0_combout ),
	.datad(av_ld_getting_data),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hFEFF;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \end_begintransfer~0 (
	.dataa(\end_begintransfer~q ),
	.datab(s0_cmd_valid),
	.datac(sink_in_reset),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\end_begintransfer~0_combout ),
	.cout());
defparam \end_begintransfer~0 .lut_mask = 16'hEFFF;
defparam \end_begintransfer~0 .sum_lutc_input = "datac";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(sink_in_reset),
	.datab(\end_begintransfer~q ),
	.datac(write_accepted1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFFFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_master_translator_1 (
	reset,
	sink_in_reset,
	waitrequest,
	mem_used_1,
	mem_used_11,
	i_read,
	read_accepted1,
	src_valid,
	uav_read,
	saved_grant_1,
	Equal2,
	saved_grant_11,
	cp_ready,
	av_readdatavalid,
	Equal1,
	take_in_data,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	sink_in_reset;
input 	waitrequest;
input 	mem_used_1;
input 	mem_used_11;
input 	i_read;
output 	read_accepted1;
input 	src_valid;
output 	uav_read;
input 	saved_grant_1;
input 	Equal2;
input 	saved_grant_11;
input 	cp_ready;
input 	av_readdatavalid;
input 	Equal1;
input 	take_in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \read_accepted~2_combout ;
wire \read_accepted~3_combout ;
wire \read_accepted~4_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb \uav_read~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read),
	.cout());
defparam \uav_read~0 .lut_mask = 16'h0FFF;
defparam \uav_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(saved_grant_11),
	.datab(waitrequest),
	.datac(mem_used_1),
	.datad(Equal1),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hBFFF;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~1 (
	.dataa(\read_accepted~0_combout ),
	.datab(saved_grant_1),
	.datac(Equal2),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFEFF;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~2 (
	.dataa(take_in_data),
	.datab(\read_accepted~1_combout ),
	.datac(src_valid),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\read_accepted~2_combout ),
	.cout());
defparam \read_accepted~2 .lut_mask = 16'hFEFF;
defparam \read_accepted~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~3 (
	.dataa(sink_in_reset),
	.datab(gnd),
	.datac(gnd),
	.datad(i_read),
	.cin(gnd),
	.combout(\read_accepted~3_combout ),
	.cout());
defparam \read_accepted~3 .lut_mask = 16'hAAFF;
defparam \read_accepted~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~4 (
	.dataa(read_accepted1),
	.datab(\read_accepted~2_combout ),
	.datac(\read_accepted~3_combout ),
	.datad(av_readdatavalid),
	.cin(gnd),
	.combout(\read_accepted~4_combout ),
	.cout());
defparam \read_accepted~4 .lut_mask = 16'hFEFF;
defparam \read_accepted~4 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_agent (
	W_alu_result_7,
	Equal3,
	always1,
	mem_used_1,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	Equal3;
input 	always1;
input 	mem_used_1;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~0 (
	.dataa(Equal3),
	.datab(always1),
	.datac(W_alu_result_7),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hEFFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_agent_1 (
	W_alu_result_24,
	Equal1,
	d_write,
	write_accepted,
	d_read,
	read_accepted,
	mem_used_128,
	Equal11,
	m0_write,
	m0_read,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_24;
input 	Equal1;
input 	d_write;
input 	write_accepted;
input 	d_read;
input 	read_accepted;
input 	mem_used_128;
input 	Equal11;
output 	m0_write;
output 	m0_read;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~2 (
	.dataa(Equal1),
	.datab(Equal11),
	.datac(W_alu_result_24),
	.datad(mem_used_128),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~2 .lut_mask = 16'hEFFF;
defparam \m0_write~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_read~2 (
	.dataa(d_read),
	.datab(read_accepted),
	.datac(m0_write),
	.datad(gnd),
	.cin(gnd),
	.combout(m0_read),
	.cout());
defparam \m0_read~2 .lut_mask = 16'hFBFB;
defparam \m0_read~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~3 (
	.dataa(d_write),
	.datab(write_accepted),
	.datac(m0_write),
	.datad(gnd),
	.cin(gnd),
	.combout(m0_write1),
	.cout());
defparam \m0_write~3 .lut_mask = 16'hFBFB;
defparam \m0_write~3 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_agent_3 (
	WideOr1,
	mem,
	local_read)/* synthesis synthesis_greybox=1 */;
input 	WideOr1;
input 	mem;
output 	local_read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \local_read~0 (
	.dataa(WideOr1),
	.datab(mem),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(local_read),
	.cout());
defparam \local_read~0 .lut_mask = 16'hEEEE;
defparam \local_read~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_agent_8 (
	mem_used_7,
	saved_grant_0,
	WideOr1,
	out_data_buffer_67,
	src_payload,
	src_payload_0,
	out_data_buffer_66,
	nonposted_write_endofpacket,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_7;
input 	saved_grant_0;
input 	WideOr1;
input 	out_data_buffer_67;
input 	src_payload;
input 	src_payload_0;
input 	out_data_buffer_66;
output 	nonposted_write_endofpacket;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \nonposted_write_endofpacket~0 (
	.dataa(WideOr1),
	.datab(src_payload),
	.datac(src_payload_0),
	.datad(out_data_buffer_66),
	.cin(gnd),
	.combout(nonposted_write_endofpacket),
	.cout());
defparam \nonposted_write_endofpacket~0 .lut_mask = 16'hFEFF;
defparam \nonposted_write_endofpacket~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~2 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_67),
	.datac(WideOr1),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~2 .lut_mask = 16'hFF7F;
defparam \m0_write~2 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_agent_9 (
	d_write,
	write_accepted,
	waitrequest_reset_override,
	saved_grant_0,
	mem_used_1,
	m0_write,
	av_waitrequest_generated,
	wait_latency_counter_1,
	cp_ready)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	waitrequest_reset_override;
input 	saved_grant_0;
input 	mem_used_1;
output 	m0_write;
input 	av_waitrequest_generated;
input 	wait_latency_counter_1;
output 	cp_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(write_accepted),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hEFFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cp_ready~0 (
	.dataa(mem_used_1),
	.datab(wait_latency_counter_1),
	.datac(waitrequest_reset_override),
	.datad(av_waitrequest_generated),
	.cin(gnd),
	.combout(cp_ready),
	.cout());
defparam \cp_ready~0 .lut_mask = 16'hEFFF;
defparam \cp_ready~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator (
	W_alu_result_7,
	Equal3,
	reset,
	read_latency_shift_reg_0,
	uav_write,
	always1,
	mem_used_1,
	wait_latency_counter_1,
	waitrequest_reset_override1,
	sink_ready,
	m0_write,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	Equal3;
input 	reset;
output 	read_latency_shift_reg_0;
input 	uav_write;
input 	always1;
input 	mem_used_1;
output 	wait_latency_counter_1;
output 	waitrequest_reset_override1;
input 	sink_ready;
input 	m0_write;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter[0]~q ;
wire \Add0~0_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter[1]~q ;
wire \wait_latency_counter[1]~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(\wait_latency_counter[1]~q ),
	.datac(Equal3),
	.datad(\wait_latency_counter[1]~0_combout ),
	.cin(gnd),
	.combout(wait_latency_counter_1),
	.cout());
defparam \wait_latency_counter[1]~1 .lut_mask = 16'hB77B;
defparam \wait_latency_counter[1]~1 .sum_lutc_input = "datac";

dffeas waitrequest_reset_override(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_reset_override1),
	.prn(vcc));
defparam waitrequest_reset_override.is_wysiwyg = "true";
defparam waitrequest_reset_override.power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(wait_latency_counter_1),
	.datac(m0_write),
	.datad(waitrequest_reset_override1),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wait_latency_counter[1]~q ),
	.datad(\wait_latency_counter[0]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(m0_write),
	.datab(waitrequest_reset_override1),
	.datac(\Add0~0_combout ),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[1]~q ),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(uav_write),
	.datab(always1),
	.datac(W_alu_result_7),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator_2 (
	reset,
	sink_in_reset,
	read_latency_shift_reg_0,
	mem_used_1,
	WideOr1,
	mem,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	sink_in_reset;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	WideOr1;
input 	mem;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(sink_in_reset),
	.datab(WideOr1),
	.datac(mem),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

endmodule

module usb_system_altera_merlin_slave_translator_3 (
	av_readdata,
	reset,
	sink_in_reset,
	read_latency_shift_reg_0,
	waitrequest,
	mem_used_1,
	local_read,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_20,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_17,
	av_readdata_pre_21,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_31,
	av_readdata_pre_30,
	av_readdata_pre_29,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	sink_in_reset;
output 	read_latency_shift_reg_0;
input 	waitrequest;
input 	mem_used_1;
input 	local_read;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_11;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	av_readdata_pre_5;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_20;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_17;
output 	av_readdata_pre_21;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_31;
output 	av_readdata_pre_30;
output 	av_readdata_pre_29;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(sink_in_reset),
	.datab(local_read),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator_4 (
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	reset,
	sink_in_reset,
	read_latency_shift_reg_0,
	uav_read,
	av_waitrequest,
	sink_ready,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	b_full,
	read_0,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_01,
	counter_reg_bit_11,
	counter_reg_bit_41,
	counter_reg_bit_51,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_22;
output 	av_readdata_pre_21;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
input 	reset;
input 	sink_in_reset;
output 	read_latency_shift_reg_0;
input 	uav_read;
input 	av_waitrequest;
input 	sink_ready;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
input 	[31:0] av_readdata;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
input 	b_full;
input 	read_0;
input 	counter_reg_bit_3;
input 	counter_reg_bit_0;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	b_full1;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_31;
input 	counter_reg_bit_21;
input 	counter_reg_bit_01;
input 	counter_reg_bit_11;
input 	counter_reg_bit_41;
input 	counter_reg_bit_51;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdata_pre[16]~7_combout ;
wire \av_readdata_pre[16]~8 ;
wire \av_readdata_pre[17]~9_combout ;
wire \av_readdata_pre[17]~10 ;
wire \av_readdata_pre[18]~11_combout ;
wire \av_readdata_pre[18]~12 ;
wire \av_readdata_pre[19]~14 ;
wire \av_readdata_pre[20]~16 ;
wire \av_readdata_pre[21]~18 ;
wire \av_readdata_pre[22]~19_combout ;
wire \av_readdata_pre[21]~17_combout ;
wire \av_readdata_pre[20]~15_combout ;
wire \av_readdata_pre[19]~13_combout ;
wire \read_latency_shift_reg~0_combout ;
wire \av_readdata_pre[13]~21_combout ;


dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(\av_readdata_pre[16]~7_combout ),
	.asdata(counter_reg_bit_01),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(\av_readdata_pre[17]~9_combout ),
	.asdata(counter_reg_bit_11),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(\av_readdata_pre[18]~11_combout ),
	.asdata(counter_reg_bit_21),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(\av_readdata_pre[22]~19_combout ),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(\av_readdata_pre[21]~17_combout ),
	.asdata(counter_reg_bit_51),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(\av_readdata_pre[20]~15_combout ),
	.asdata(counter_reg_bit_41),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(\av_readdata_pre[19]~13_combout ),
	.asdata(counter_reg_bit_31),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

cycloneive_lcell_comb \av_readdata_pre[16]~7 (
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\av_readdata_pre[16]~7_combout ),
	.cout(\av_readdata_pre[16]~8 ));
defparam \av_readdata_pre[16]~7 .lut_mask = 16'hAA55;
defparam \av_readdata_pre[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[17]~9 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[16]~8 ),
	.combout(\av_readdata_pre[17]~9_combout ),
	.cout(\av_readdata_pre[17]~10 ));
defparam \av_readdata_pre[17]~9 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[17]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[18]~11 (
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[17]~10 ),
	.combout(\av_readdata_pre[18]~11_combout ),
	.cout(\av_readdata_pre[18]~12 ));
defparam \av_readdata_pre[18]~11 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[18]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[19]~13 (
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[18]~12 ),
	.combout(\av_readdata_pre[19]~13_combout ),
	.cout(\av_readdata_pre[19]~14 ));
defparam \av_readdata_pre[19]~13 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[19]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[20]~15 (
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[19]~14 ),
	.combout(\av_readdata_pre[20]~15_combout ),
	.cout(\av_readdata_pre[20]~16 ));
defparam \av_readdata_pre[20]~15 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[20]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[21]~17 (
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[20]~16 ),
	.combout(\av_readdata_pre[21]~17_combout ),
	.cout(\av_readdata_pre[21]~18 ));
defparam \av_readdata_pre[21]~17 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[21]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[22]~19 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\av_readdata_pre[21]~18 ),
	.combout(\av_readdata_pre[22]~19_combout ),
	.cout());
defparam \av_readdata_pre[22]~19 .lut_mask = 16'h5A5A;
defparam \av_readdata_pre[22]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(sink_in_reset),
	.datab(uav_read),
	.datac(av_waitrequest),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[13]~21 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_readdata_pre[13]~21_combout ),
	.cout());
defparam \av_readdata_pre[13]~21 .lut_mask = 16'h5555;
defparam \av_readdata_pre[13]~21 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator_5 (
	W_alu_result_7,
	W_alu_result_4,
	W_alu_result_5,
	reset,
	Equal3,
	mem_used_1,
	always0,
	d_write,
	write_accepted,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg,
	sink_in_reset,
	d_read,
	read_accepted,
	read_latency_shift_reg1,
	read_latency_shift_reg_0,
	uav_write,
	s0_cmd_valid,
	Equal6,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	reset;
input 	Equal3;
input 	mem_used_1;
input 	always0;
input 	d_write;
input 	write_accepted;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg;
input 	sink_in_reset;
input 	d_read;
input 	read_accepted;
output 	read_latency_shift_reg1;
output 	read_latency_shift_reg_0;
input 	uav_write;
input 	s0_cmd_valid;
input 	Equal6;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter[1]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \read_latency_shift_reg~0_combout ;
wire \read_latency_shift_reg~1_combout ;
wire \read_latency_shift_reg~4_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(wait_latency_counter_1),
	.datab(Equal3),
	.datac(\read_latency_shift_reg~0_combout ),
	.datad(\read_latency_shift_reg~1_combout ),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hFFFD;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~3 (
	.dataa(sink_in_reset),
	.datab(d_read),
	.datac(gnd),
	.datad(read_accepted),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~3 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~3 .sum_lutc_input = "datac";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(wait_latency_counter_0),
	.datab(always0),
	.datac(uav_write),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'h96FF;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(always0),
	.datab(sink_in_reset),
	.datac(s0_cmd_valid),
	.datad(\wait_latency_counter[1]~0_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~1_combout ),
	.cout());
defparam \wait_latency_counter[1]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[1]~1_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[1]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(wait_latency_counter_0),
	.datab(d_write),
	.datac(mem_used_1),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'h6996;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(W_alu_result_7),
	.datab(W_alu_result_4),
	.datac(W_alu_result_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hBFBF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~4 (
	.dataa(Equal6),
	.datab(\wait_latency_counter[1]~0_combout ),
	.datac(read_latency_shift_reg1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~4_combout ),
	.cout());
defparam \read_latency_shift_reg~4 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~4 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator_6 (
	W_alu_result_4,
	W_alu_result_5,
	reset,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	uav_write,
	waitrequest_reset_override,
	uav_read,
	always1,
	wait_latency_counter_01,
	s0_cmd_valid,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	reset;
input 	mem_used_1;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
input 	uav_write;
input 	waitrequest_reset_override;
input 	uav_read;
input 	always1;
output 	wait_latency_counter_01;
input 	s0_cmd_valid;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter~4_combout ;
wire \wait_latency_counter[0]~0_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(wait_latency_counter_0),
	.datab(wait_latency_counter_1),
	.datac(always1),
	.datad(\wait_latency_counter[0]~0_combout ),
	.cin(gnd),
	.combout(wait_latency_counter_01),
	.cout());
defparam \wait_latency_counter[0]~1 .lut_mask = 16'hB77B;
defparam \wait_latency_counter[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(always0),
	.datab(uav_read),
	.datac(waitrequest_reset_override),
	.datad(wait_latency_counter_01),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~2 (
	.dataa(always0),
	.datab(waitrequest_reset_override),
	.datac(s0_cmd_valid),
	.datad(wait_latency_counter_01),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~2_combout ),
	.cout());
defparam \wait_latency_counter[0]~2 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[0]~2_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~4 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[0]~2_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~4_combout ),
	.cout());
defparam \wait_latency_counter~4 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(uav_write),
	.datab(W_alu_result_4),
	.datac(W_alu_result_5),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'hFF7F;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator_7 (
	W_alu_result_4,
	W_alu_result_5,
	reset,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	uav_write,
	waitrequest_reset_override,
	uav_read,
	always1,
	wait_latency_counter_11,
	s0_cmd_valid,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	reset;
input 	mem_used_1;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
input 	uav_write;
input 	waitrequest_reset_override;
input 	uav_read;
input 	always1;
output 	wait_latency_counter_11;
input 	s0_cmd_valid;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~2_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter~4_combout ;
wire \wait_latency_counter[1]~0_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(wait_latency_counter_0),
	.datab(wait_latency_counter_1),
	.datac(always1),
	.datad(\wait_latency_counter[1]~0_combout ),
	.cin(gnd),
	.combout(wait_latency_counter_11),
	.cout());
defparam \wait_latency_counter[1]~1 .lut_mask = 16'hB77B;
defparam \wait_latency_counter[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(always0),
	.datab(uav_read),
	.datac(waitrequest_reset_override),
	.datad(wait_latency_counter_11),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~2 (
	.dataa(always0),
	.datab(waitrequest_reset_override),
	.datac(s0_cmd_valid),
	.datad(wait_latency_counter_11),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~2_combout ),
	.cout());
defparam \wait_latency_counter[1]~2 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[1]~2_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~4 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[1]~2_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~4_combout ),
	.cout());
defparam \wait_latency_counter~4 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(uav_write),
	.datab(W_alu_result_4),
	.datac(W_alu_result_5),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_slave_translator_9 (
	reset,
	read_latency_shift_reg_0,
	waitrequest_reset_override,
	sink_ready,
	saved_grant_1,
	src_valid,
	mem_used_1,
	m0_write,
	av_waitrequest_generated,
	wait_latency_counter_1,
	src_data_68,
	always1,
	read_latency_shift_reg,
	WideOr1,
	src_payload,
	av_readdata_pre_30,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	read_latency_shift_reg_0;
input 	waitrequest_reset_override;
input 	sink_ready;
input 	saved_grant_1;
input 	src_valid;
input 	mem_used_1;
input 	m0_write;
output 	av_waitrequest_generated;
output 	wait_latency_counter_1;
input 	src_data_68;
input 	always1;
output 	read_latency_shift_reg;
input 	WideOr1;
input 	src_payload;
output 	av_readdata_pre_30;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~2_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~3_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \av_waitrequest_generated~0 (
	.dataa(sink_ready),
	.datab(src_valid),
	.datac(\wait_latency_counter[0]~q ),
	.datad(m0_write),
	.cin(gnd),
	.combout(av_waitrequest_generated),
	.cout());
defparam \av_waitrequest_generated~0 .lut_mask = 16'h6996;
defparam \av_waitrequest_generated~0 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(waitrequest_reset_override),
	.datab(av_waitrequest_generated),
	.datac(\read_latency_shift_reg~0_combout ),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(read_latency_shift_reg),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~2_combout ),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hAAFF;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(waitrequest_reset_override),
	.datab(src_payload),
	.datac(src_data_68),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(WideOr1),
	.datab(\wait_latency_counter[0]~0_combout ),
	.datac(wait_latency_counter_1),
	.datad(av_waitrequest_generated),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.cout());
defparam \wait_latency_counter[0]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[0]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[0]~1_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(\wait_latency_counter[0]~q ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(src_data_68),
	.datab(sink_ready),
	.datac(saved_grant_1),
	.datad(always1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_cmd_demux (
	W_alu_result_7,
	W_alu_result_4,
	W_alu_result_5,
	Equal3,
	mem_used_1,
	always0,
	always01,
	read_latency_shift_reg,
	sink_in_reset,
	Equal2,
	saved_grant_0,
	waitrequest,
	mem_used_11,
	always1,
	mem_used_12,
	wait_latency_counter_1,
	waitrequest_reset_override,
	saved_grant_01,
	mem_used_13,
	full,
	mem_used_128,
	Equal1,
	saved_grant_02,
	always11,
	sink_ready,
	mem_used_14,
	av_waitrequest_generated,
	wait_latency_counter_11,
	mem_used_15,
	Equal9,
	av_waitrequest,
	sink_ready1,
	in_data_toggle,
	dreg_0,
	Equal91,
	wait_latency_counter_12,
	wait_latency_counter_0,
	WideOr0,
	sink_ready2,
	always12,
	sink_ready3,
	sink_ready4,
	always13,
	sink_ready5)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	Equal3;
input 	mem_used_1;
input 	always0;
input 	always01;
input 	read_latency_shift_reg;
input 	sink_in_reset;
input 	Equal2;
input 	saved_grant_0;
input 	waitrequest;
input 	mem_used_11;
input 	always1;
input 	mem_used_12;
input 	wait_latency_counter_1;
input 	waitrequest_reset_override;
input 	saved_grant_01;
input 	mem_used_13;
input 	full;
input 	mem_used_128;
input 	Equal1;
input 	saved_grant_02;
input 	always11;
output 	sink_ready;
input 	mem_used_14;
input 	av_waitrequest_generated;
input 	wait_latency_counter_11;
input 	mem_used_15;
input 	Equal9;
input 	av_waitrequest;
output 	sink_ready1;
input 	in_data_toggle;
input 	dreg_0;
input 	Equal91;
input 	wait_latency_counter_12;
input 	wait_latency_counter_0;
output 	WideOr0;
output 	sink_ready2;
input 	always12;
output 	sink_ready3;
output 	sink_ready4;
input 	always13;
output 	sink_ready5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \sink_ready~1_combout ;
wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \WideOr0~2_combout ;
wire \WideOr0~3_combout ;
wire \WideOr0~4_combout ;
wire \sink_ready~3_combout ;
wire \sink_ready~4_combout ;
wire \sink_ready~5_combout ;
wire \sink_ready~6_combout ;
wire \sink_ready~8_combout ;
wire \sink_ready~9_combout ;
wire \sink_ready~10_combout ;
wire \WideOr0~5_combout ;
wire \WideOr0~6_combout ;


cycloneive_lcell_comb \sink_ready~2 (
	.dataa(W_alu_result_7),
	.datab(Equal3),
	.datac(saved_grant_02),
	.datad(always11),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~2 .lut_mask = 16'hFFFE;
defparam \sink_ready~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~7 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_7),
	.datac(W_alu_result_4),
	.datad(Equal3),
	.cin(gnd),
	.combout(sink_ready1),
	.cout());
defparam \sink_ready~7 .lut_mask = 16'h8BFF;
defparam \sink_ready~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~7 (
	.dataa(\WideOr0~0_combout ),
	.datab(\WideOr0~4_combout ),
	.datac(\sink_ready~4_combout ),
	.datad(\WideOr0~6_combout ),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~7 .lut_mask = 16'hFFFE;
defparam \WideOr0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~11 (
	.dataa(W_alu_result_7),
	.datab(Equal3),
	.datac(Equal9),
	.datad(mem_used_15),
	.cin(gnd),
	.combout(sink_ready2),
	.cout());
defparam \sink_ready~11 .lut_mask = 16'hFEFF;
defparam \sink_ready~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~12 (
	.dataa(always12),
	.datab(wait_latency_counter_1),
	.datac(waitrequest_reset_override),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(sink_ready3),
	.cout());
defparam \sink_ready~12 .lut_mask = 16'hFEFF;
defparam \sink_ready~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~13 (
	.dataa(always12),
	.datab(wait_latency_counter_1),
	.datac(waitrequest_reset_override),
	.datad(gnd),
	.cin(gnd),
	.combout(sink_ready4),
	.cout());
defparam \sink_ready~13 .lut_mask = 16'hFEFE;
defparam \sink_ready~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~14 (
	.dataa(\sink_ready~9_combout ),
	.datab(always12),
	.datac(always13),
	.datad(Equal91),
	.cin(gnd),
	.combout(sink_ready5),
	.cout());
defparam \sink_ready~14 .lut_mask = 16'hBFFF;
defparam \sink_ready~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~0 (
	.dataa(Equal2),
	.datab(saved_grant_0),
	.datac(waitrequest),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(\sink_ready~0_combout ),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hEFFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~1 (
	.dataa(Equal3),
	.datab(always1),
	.datac(waitrequest_reset_override),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(\sink_ready~1_combout ),
	.cout());
defparam \sink_ready~1 .lut_mask = 16'hFEFF;
defparam \sink_ready~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\sink_ready~0_combout ),
	.datab(wait_latency_counter_1),
	.datac(\sink_ready~1_combout ),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hFEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~1 (
	.dataa(mem_used_13),
	.datab(W_alu_result_4),
	.datac(W_alu_result_7),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(\WideOr0~1_combout ),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hFDFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~2 (
	.dataa(full),
	.datab(mem_used_128),
	.datac(Equal1),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr0~2_combout ),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'h7F7F;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~3 (
	.dataa(saved_grant_01),
	.datab(Equal3),
	.datac(\WideOr0~1_combout ),
	.datad(\WideOr0~2_combout ),
	.cin(gnd),
	.combout(\WideOr0~3_combout ),
	.cout());
defparam \WideOr0~3 .lut_mask = 16'hFFFE;
defparam \WideOr0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~4 (
	.dataa(sink_in_reset),
	.datab(\WideOr0~3_combout ),
	.datac(read_latency_shift_reg),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\WideOr0~4_combout ),
	.cout());
defparam \WideOr0~4 .lut_mask = 16'hFEFF;
defparam \WideOr0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~3 (
	.dataa(mem_used_14),
	.datab(wait_latency_counter_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_ready~3_combout ),
	.cout());
defparam \sink_ready~3 .lut_mask = 16'h7777;
defparam \sink_ready~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~4 (
	.dataa(sink_ready),
	.datab(waitrequest_reset_override),
	.datac(av_waitrequest_generated),
	.datad(\sink_ready~3_combout ),
	.cin(gnd),
	.combout(\sink_ready~4_combout ),
	.cout());
defparam \sink_ready~4 .lut_mask = 16'hFFFE;
defparam \sink_ready~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~5 (
	.dataa(av_waitrequest),
	.datab(W_alu_result_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_ready~5_combout ),
	.cout());
defparam \sink_ready~5 .lut_mask = 16'hEEEE;
defparam \sink_ready~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~6 (
	.dataa(mem_used_15),
	.datab(Equal3),
	.datac(Equal9),
	.datad(\sink_ready~5_combout ),
	.cin(gnd),
	.combout(\sink_ready~6_combout ),
	.cout());
defparam \sink_ready~6 .lut_mask = 16'hFFFD;
defparam \sink_ready~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~8 (
	.dataa(W_alu_result_7),
	.datab(always1),
	.datac(always11),
	.datad(Equal3),
	.cin(gnd),
	.combout(\sink_ready~8_combout ),
	.cout());
defparam \sink_ready~8 .lut_mask = 16'h27FF;
defparam \sink_ready~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~9 (
	.dataa(Equal1),
	.datab(in_data_toggle),
	.datac(dreg_0),
	.datad(Equal2),
	.cin(gnd),
	.combout(\sink_ready~9_combout ),
	.cout());
defparam \sink_ready~9 .lut_mask = 16'hBEFF;
defparam \sink_ready~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~10 (
	.dataa(sink_ready1),
	.datab(\sink_ready~8_combout ),
	.datac(\sink_ready~9_combout ),
	.datad(Equal91),
	.cin(gnd),
	.combout(\sink_ready~10_combout ),
	.cout());
defparam \sink_ready~10 .lut_mask = 16'hFEFF;
defparam \sink_ready~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~5 (
	.dataa(always0),
	.datab(always01),
	.datac(wait_latency_counter_12),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\WideOr0~5_combout ),
	.cout());
defparam \WideOr0~5 .lut_mask = 16'hFFFE;
defparam \WideOr0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~6 (
	.dataa(\sink_ready~6_combout ),
	.datab(\sink_ready~10_combout ),
	.datac(waitrequest_reset_override),
	.datad(\WideOr0~5_combout ),
	.cin(gnd),
	.combout(\WideOr0~6_combout ),
	.cout());
defparam \WideOr0~6 .lut_mask = 16'hFFFE;
defparam \WideOr0~6 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_cmd_demux_001 (
	Equal1,
	F_pc_10,
	F_pc_9,
	i_read,
	read_accepted,
	uav_read,
	Equal2,
	src1_valid,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	Equal1;
input 	F_pc_10;
input 	F_pc_9;
input 	i_read;
input 	read_accepted;
input 	uav_read;
input 	Equal2;
output 	src1_valid;
output 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src1_valid~0 (
	.dataa(Equal1),
	.datab(F_pc_9),
	.datac(uav_read),
	.datad(F_pc_10),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFF;
defparam \src1_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src2_valid~0 (
	.dataa(Equal2),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted),
	.cin(gnd),
	.combout(src2_valid),
	.cout());
defparam \src2_valid~0 .lut_mask = 16'hAFFF;
defparam \src2_valid~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_cmd_mux_001 (
	W_alu_result_2,
	Equal6,
	d_write,
	write_accepted,
	altera_reset_synchronizer_int_chain_out,
	saved_grant_0,
	uav_read,
	always1,
	saved_grant_1,
	Equal1,
	Equal2,
	always11,
	src_valid,
	uav_read1,
	F_pc_0,
	src_data_68,
	always12,
	always13,
	WideOr11,
	cp_ready,
	src_payload,
	src_data_38,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
input 	Equal6;
input 	d_write;
input 	write_accepted;
input 	altera_reset_synchronizer_int_chain_out;
output 	saved_grant_0;
input 	uav_read;
input 	always1;
output 	saved_grant_1;
input 	Equal1;
input 	Equal2;
input 	always11;
output 	src_valid;
input 	uav_read1;
input 	F_pc_0;
output 	src_data_68;
input 	always12;
input 	always13;
output 	WideOr11;
input 	cp_ready;
output 	src_payload;
output 	src_data_38;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;


usb_system_altera_merlin_arbitrator arb(
	.reset(altera_reset_synchronizer_int_chain_out),
	.always1(always12),
	.always11(always13),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.WideOr1(WideOr11),
	.packet_in_progress(\packet_in_progress~q ),
	.cp_ready(cp_ready),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(saved_grant_1),
	.datab(Equal1),
	.datac(Equal2),
	.datad(always11),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hFFFE;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[68] (
	.dataa(uav_read),
	.datab(saved_grant_1),
	.datac(uav_read1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_68),
	.cout());
defparam \src_data[68] .lut_mask = 16'hFFFE;
defparam \src_data[68] .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(src_valid),
	.datab(Equal6),
	.datac(saved_grant_0),
	.datad(always1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(saved_grant_1),
	.datac(F_pc_0),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEEEE;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(\packet_in_progress~q ),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h8BFF;
defparam \update_grant~1 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_arbitrator (
	reset,
	always1,
	always11,
	grant_0,
	update_grant,
	WideOr1,
	packet_in_progress,
	cp_ready,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	always1;
input 	always11;
output 	grant_0;
input 	update_grant;
input 	WideOr1;
input 	packet_in_progress;
input 	cp_ready;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(always11),
	.datab(\top_priority_reg[1]~q ),
	.datac(always1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(always1),
	.datab(\top_priority_reg[1]~q ),
	.datac(always11),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(WideOr1),
	.datac(packet_in_progress),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hF7D5;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(always11),
	.datab(always1),
	.datac(\top_priority_reg[0]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'hEFEF;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~2 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.cout());
defparam \top_priority_reg[0]~2 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~2 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module usb_system_usb_system_mm_interconnect_0_cmd_mux_001_1 (
	W_alu_result_7,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_6,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	Equal2,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	F_pc_8,
	F_pc_7,
	F_pc_5,
	F_pc_6,
	F_pc_4,
	F_pc_1,
	F_pc_3,
	F_pc_2,
	s0_cmd_valid,
	F_pc_0,
	src1_valid,
	saved_grant_1,
	WideOr11,
	hbreak_enabled,
	src_data_46,
	d_byteenable_0,
	d_byteenable_1,
	d_byteenable_2,
	d_byteenable_3,
	src_payload,
	src_payload1,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_22,
	d_writedata_23,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_34,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_35,
	src_payload12,
	src_payload13,
	src_payload14,
	src_data_33,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_6;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	Equal2;
output 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_4;
input 	F_pc_1;
input 	F_pc_3;
input 	F_pc_2;
input 	s0_cmd_valid;
input 	F_pc_0;
input 	src1_valid;
output 	saved_grant_1;
output 	WideOr11;
input 	hbreak_enabled;
output 	src_data_46;
input 	d_byteenable_0;
input 	d_byteenable_1;
input 	d_byteenable_2;
input 	d_byteenable_3;
output 	src_payload;
output 	src_payload1;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_22;
input 	d_writedata_23;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_data_34;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_data_35;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_data_33;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~0_combout ;


usb_system_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.Equal2(Equal2),
	.s0_cmd_valid(s0_cmd_valid),
	.src1_valid(src1_valid),
	.src_valid(\src_valid~0_combout ),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(src1_valid),
	.datac(saved_grant_1),
	.datad(\src_valid~0_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(W_alu_result_10),
	.datab(F_pc_8),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(W_alu_result_4),
	.datab(F_pc_2),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(W_alu_result_5),
	.datab(F_pc_3),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(W_alu_result_6),
	.datab(F_pc_4),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(W_alu_result_7),
	.datab(F_pc_5),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(W_alu_result_8),
	.datab(F_pc_6),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(W_alu_result_9),
	.datab(F_pc_7),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(d_writedata_11),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(d_writedata_13),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(d_writedata_16),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(d_writedata_12),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(d_writedata_14),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(d_writedata_15),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(d_writedata_10),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(d_writedata_9),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(d_writedata_8),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(d_writedata_17),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEFFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(Equal2),
	.datab(s0_cmd_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hEEEE;
defparam \src_valid~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_arbitrator_1 (
	reset,
	Equal2,
	s0_cmd_valid,
	src1_valid,
	src_valid,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	Equal2;
input 	s0_cmd_valid;
input 	src1_valid;
input 	src_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~3_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src1_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src1_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(\top_priority_reg[0]~q ),
	.datad(src_valid),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~2 (
	.dataa(Equal2),
	.datab(s0_cmd_valid),
	.datac(update_grant),
	.datad(src1_valid),
	.cin(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.cout());
defparam \top_priority_reg[0]~2 .lut_mask = 16'hFFFE;
defparam \top_priority_reg[0]~2 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~2_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~3 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~3_combout ),
	.cout());
defparam \top_priority_reg[0]~3 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~3 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~2_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module usb_system_usb_system_mm_interconnect_0_cmd_mux_001_2 (
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	r_sync_rst,
	Equal6,
	sink_in_reset,
	saved_grant_0,
	mem_used_1,
	F_pc_1,
	i_read,
	read_accepted,
	s0_cmd_valid,
	saved_grant_1,
	Equal2,
	Equal7,
	WideOr11,
	F_pc_0,
	src_data_38,
	src_data_39,
	src2_valid,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	r_sync_rst;
input 	Equal6;
input 	sink_in_reset;
output 	saved_grant_0;
input 	mem_used_1;
input 	F_pc_1;
input 	i_read;
input 	read_accepted;
input 	s0_cmd_valid;
output 	saved_grant_1;
input 	Equal2;
input 	Equal7;
output 	WideOr11;
input 	F_pc_0;
output 	src_data_38;
output 	src_data_39;
input 	src2_valid;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_valid~2_combout ;
wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~3_combout ;


usb_system_altera_merlin_arbitrator_2 arb(
	.reset(r_sync_rst),
	.src_valid(\src_valid~2_combout ),
	.src2_valid(src2_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

cycloneive_lcell_comb \src_valid~2 (
	.dataa(W_alu_result_4),
	.datab(Equal6),
	.datac(s0_cmd_valid),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(\src_valid~2_combout ),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hFEFF;
defparam \src_valid~2 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(\src_valid~3_combout ),
	.datab(Equal7),
	.datac(saved_grant_0),
	.datad(s0_cmd_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(saved_grant_1),
	.datac(F_pc_0),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(sink_in_reset),
	.datab(saved_grant_0),
	.datac(saved_grant_1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFEFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~3 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(saved_grant_1),
	.datad(Equal2),
	.cin(gnd),
	.combout(\src_valid~3_combout ),
	.cout());
defparam \src_valid~3 .lut_mask = 16'hFFF7;
defparam \src_valid~3 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_arbitrator_2 (
	reset,
	src_valid,
	src2_valid,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src_valid;
input 	src2_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src2_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src2_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src2_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module usb_system_usb_system_mm_interconnect_0_cmd_mux_001_3 (
	wire_pll7_clk_0,
	entries_1,
	entries_0,
	altera_reset_synchronizer_int_chain_out,
	mem_used_7,
	last_cycle,
	saved_grant_0,
	saved_grant_1,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	WideOr11,
	out_data_buffer_67,
	src_payload,
	out_data_buffer_68,
	out_data_buffer_681,
	src_data_68,
	out_data_buffer_48,
	out_data_buffer_481,
	src_data_48,
	out_data_buffer_62,
	out_data_buffer_621,
	src_data_62,
	out_data_buffer_49,
	out_data_buffer_491,
	src_data_49,
	out_data_buffer_51,
	out_data_buffer_511,
	src_data_51,
	out_data_buffer_50,
	out_data_buffer_501,
	src_data_50,
	out_data_buffer_53,
	out_data_buffer_531,
	src_data_53,
	out_data_buffer_52,
	out_data_buffer_521,
	src_data_52,
	out_data_buffer_55,
	out_data_buffer_551,
	src_data_55,
	out_data_buffer_54,
	out_data_buffer_541,
	src_data_54,
	out_data_buffer_57,
	out_data_buffer_571,
	src_data_57,
	out_data_buffer_56,
	out_data_buffer_561,
	src_data_56,
	out_data_buffer_59,
	out_data_buffer_591,
	src_data_59,
	out_data_buffer_58,
	out_data_buffer_581,
	src_data_58,
	out_data_buffer_61,
	out_data_buffer_611,
	src_data_61,
	out_data_buffer_60,
	out_data_buffer_601,
	src_data_60,
	out_data_buffer_38,
	out_data_buffer_381,
	src_data_38,
	out_data_buffer_39,
	out_data_buffer_391,
	src_data_39,
	out_data_buffer_40,
	out_data_buffer_401,
	src_data_40,
	out_data_buffer_41,
	out_data_buffer_411,
	src_data_41,
	out_data_buffer_42,
	out_data_buffer_421,
	src_data_42,
	out_data_buffer_43,
	out_data_buffer_431,
	src_data_43,
	out_data_buffer_44,
	out_data_buffer_441,
	src_data_44,
	out_data_buffer_45,
	out_data_buffer_451,
	src_data_45,
	out_data_buffer_46,
	out_data_buffer_461,
	src_data_46,
	out_data_buffer_47,
	out_data_buffer_471,
	src_data_47,
	out_data_buffer_107,
	out_data_buffer_1071,
	src_payload_0,
	out_data_buffer_0,
	src_payload1,
	out_data_buffer_1,
	src_payload2,
	out_data_buffer_2,
	src_payload3,
	out_data_buffer_3,
	src_payload4,
	out_data_buffer_4,
	src_payload5,
	out_data_buffer_5,
	src_payload6,
	out_data_buffer_6,
	src_payload7,
	out_data_buffer_7,
	src_payload8,
	out_data_buffer_8,
	src_payload9,
	out_data_buffer_9,
	src_payload10,
	out_data_buffer_10,
	src_payload11,
	out_data_buffer_11,
	src_payload12,
	out_data_buffer_12,
	src_payload13,
	out_data_buffer_13,
	src_payload14,
	out_data_buffer_14,
	src_payload15,
	out_data_buffer_15,
	src_payload16,
	out_data_buffer_16,
	src_payload17,
	out_data_buffer_17,
	src_payload18,
	out_data_buffer_18,
	src_payload19,
	out_data_buffer_19,
	src_payload20,
	out_data_buffer_20,
	src_payload21,
	out_data_buffer_21,
	src_payload22,
	out_data_buffer_22,
	src_payload23,
	out_data_buffer_23,
	src_payload24,
	out_data_buffer_24,
	src_payload25,
	out_data_buffer_25,
	src_payload26,
	out_data_buffer_26,
	src_payload27,
	out_data_buffer_27,
	src_payload28,
	out_data_buffer_28,
	src_payload29,
	out_data_buffer_29,
	src_payload30,
	out_data_buffer_30,
	src_payload31,
	out_data_buffer_31,
	src_payload32)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	entries_1;
input 	entries_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	mem_used_7;
output 	last_cycle;
output 	saved_grant_0;
output 	saved_grant_1;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
output 	WideOr11;
input 	out_data_buffer_67;
output 	src_payload;
input 	out_data_buffer_68;
input 	out_data_buffer_681;
output 	src_data_68;
input 	out_data_buffer_48;
input 	out_data_buffer_481;
output 	src_data_48;
input 	out_data_buffer_62;
input 	out_data_buffer_621;
output 	src_data_62;
input 	out_data_buffer_49;
input 	out_data_buffer_491;
output 	src_data_49;
input 	out_data_buffer_51;
input 	out_data_buffer_511;
output 	src_data_51;
input 	out_data_buffer_50;
input 	out_data_buffer_501;
output 	src_data_50;
input 	out_data_buffer_53;
input 	out_data_buffer_531;
output 	src_data_53;
input 	out_data_buffer_52;
input 	out_data_buffer_521;
output 	src_data_52;
input 	out_data_buffer_55;
input 	out_data_buffer_551;
output 	src_data_55;
input 	out_data_buffer_54;
input 	out_data_buffer_541;
output 	src_data_54;
input 	out_data_buffer_57;
input 	out_data_buffer_571;
output 	src_data_57;
input 	out_data_buffer_56;
input 	out_data_buffer_561;
output 	src_data_56;
input 	out_data_buffer_59;
input 	out_data_buffer_591;
output 	src_data_59;
input 	out_data_buffer_58;
input 	out_data_buffer_581;
output 	src_data_58;
input 	out_data_buffer_61;
input 	out_data_buffer_611;
output 	src_data_61;
input 	out_data_buffer_60;
input 	out_data_buffer_601;
output 	src_data_60;
input 	out_data_buffer_38;
input 	out_data_buffer_381;
output 	src_data_38;
input 	out_data_buffer_39;
input 	out_data_buffer_391;
output 	src_data_39;
input 	out_data_buffer_40;
input 	out_data_buffer_401;
output 	src_data_40;
input 	out_data_buffer_41;
input 	out_data_buffer_411;
output 	src_data_41;
input 	out_data_buffer_42;
input 	out_data_buffer_421;
output 	src_data_42;
input 	out_data_buffer_43;
input 	out_data_buffer_431;
output 	src_data_43;
input 	out_data_buffer_44;
input 	out_data_buffer_441;
output 	src_data_44;
input 	out_data_buffer_45;
input 	out_data_buffer_451;
output 	src_data_45;
input 	out_data_buffer_46;
input 	out_data_buffer_461;
output 	src_data_46;
input 	out_data_buffer_47;
input 	out_data_buffer_471;
output 	src_data_47;
input 	out_data_buffer_107;
input 	out_data_buffer_1071;
output 	src_payload_0;
input 	out_data_buffer_0;
output 	src_payload1;
input 	out_data_buffer_1;
output 	src_payload2;
input 	out_data_buffer_2;
output 	src_payload3;
input 	out_data_buffer_3;
output 	src_payload4;
input 	out_data_buffer_4;
output 	src_payload5;
input 	out_data_buffer_5;
output 	src_payload6;
input 	out_data_buffer_6;
output 	src_payload7;
input 	out_data_buffer_7;
output 	src_payload8;
input 	out_data_buffer_8;
output 	src_payload9;
input 	out_data_buffer_9;
output 	src_payload10;
input 	out_data_buffer_10;
output 	src_payload11;
input 	out_data_buffer_11;
output 	src_payload12;
input 	out_data_buffer_12;
output 	src_payload13;
input 	out_data_buffer_13;
output 	src_payload14;
input 	out_data_buffer_14;
output 	src_payload15;
input 	out_data_buffer_15;
output 	src_payload16;
input 	out_data_buffer_16;
output 	src_payload17;
input 	out_data_buffer_17;
output 	src_payload18;
input 	out_data_buffer_18;
output 	src_payload19;
input 	out_data_buffer_19;
output 	src_payload20;
input 	out_data_buffer_20;
output 	src_payload21;
input 	out_data_buffer_21;
output 	src_payload22;
input 	out_data_buffer_22;
output 	src_payload23;
input 	out_data_buffer_23;
output 	src_payload24;
input 	out_data_buffer_24;
output 	src_payload25;
input 	out_data_buffer_25;
output 	src_payload26;
input 	out_data_buffer_26;
output 	src_payload27;
input 	out_data_buffer_27;
output 	src_payload28;
input 	out_data_buffer_28;
output 	src_payload29;
input 	out_data_buffer_29;
output 	src_payload30;
input 	out_data_buffer_30;
output 	src_payload31;
input 	out_data_buffer_31;
output 	src_payload32;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


usb_system_altera_merlin_arbitrator_3 arb(
	.clk(wire_pll7_clk_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid1),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.grant_1(\arb|grant[1]~1_combout ));

cycloneive_lcell_comb \last_cycle~0 (
	.dataa(entries_0),
	.datab(gnd),
	.datac(entries_1),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(last_cycle),
	.cout());
defparam \last_cycle~0 .lut_mask = 16'hAFFF;
defparam \last_cycle~0 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_valid),
	.datad(out_valid1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_67),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[68] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_68),
	.datad(out_data_buffer_681),
	.cin(gnd),
	.combout(src_data_68),
	.cout());
defparam \src_data[68] .lut_mask = 16'hFFFE;
defparam \src_data[68] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[48] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_48),
	.datad(out_data_buffer_481),
	.cin(gnd),
	.combout(src_data_48),
	.cout());
defparam \src_data[48] .lut_mask = 16'hFFFE;
defparam \src_data[48] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[62] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_62),
	.datad(out_data_buffer_621),
	.cin(gnd),
	.combout(src_data_62),
	.cout());
defparam \src_data[62] .lut_mask = 16'hFFFE;
defparam \src_data[62] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[49] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_49),
	.datad(out_data_buffer_491),
	.cin(gnd),
	.combout(src_data_49),
	.cout());
defparam \src_data[49] .lut_mask = 16'hFFFE;
defparam \src_data[49] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[51] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_51),
	.datad(out_data_buffer_511),
	.cin(gnd),
	.combout(src_data_51),
	.cout());
defparam \src_data[51] .lut_mask = 16'hFFFE;
defparam \src_data[51] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[50] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_50),
	.datad(out_data_buffer_501),
	.cin(gnd),
	.combout(src_data_50),
	.cout());
defparam \src_data[50] .lut_mask = 16'hFFFE;
defparam \src_data[50] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[53] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_53),
	.datad(out_data_buffer_531),
	.cin(gnd),
	.combout(src_data_53),
	.cout());
defparam \src_data[53] .lut_mask = 16'hFFFE;
defparam \src_data[53] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[52] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_52),
	.datad(out_data_buffer_521),
	.cin(gnd),
	.combout(src_data_52),
	.cout());
defparam \src_data[52] .lut_mask = 16'hFFFE;
defparam \src_data[52] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[55] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_55),
	.datad(out_data_buffer_551),
	.cin(gnd),
	.combout(src_data_55),
	.cout());
defparam \src_data[55] .lut_mask = 16'hFFFE;
defparam \src_data[55] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[54] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_54),
	.datad(out_data_buffer_541),
	.cin(gnd),
	.combout(src_data_54),
	.cout());
defparam \src_data[54] .lut_mask = 16'hFFFE;
defparam \src_data[54] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[57] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_57),
	.datad(out_data_buffer_571),
	.cin(gnd),
	.combout(src_data_57),
	.cout());
defparam \src_data[57] .lut_mask = 16'hFFFE;
defparam \src_data[57] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[56] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_56),
	.datad(out_data_buffer_561),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[59] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_59),
	.datad(out_data_buffer_591),
	.cin(gnd),
	.combout(src_data_59),
	.cout());
defparam \src_data[59] .lut_mask = 16'hFFFE;
defparam \src_data[59] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[58] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_58),
	.datad(out_data_buffer_581),
	.cin(gnd),
	.combout(src_data_58),
	.cout());
defparam \src_data[58] .lut_mask = 16'hFFFE;
defparam \src_data[58] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[61] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_61),
	.datad(out_data_buffer_611),
	.cin(gnd),
	.combout(src_data_61),
	.cout());
defparam \src_data[61] .lut_mask = 16'hFFFE;
defparam \src_data[61] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[60] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_60),
	.datad(out_data_buffer_601),
	.cin(gnd),
	.combout(src_data_60),
	.cout());
defparam \src_data[60] .lut_mask = 16'hFFFE;
defparam \src_data[60] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_38),
	.datad(out_data_buffer_381),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_39),
	.datad(out_data_buffer_391),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_40),
	.datad(out_data_buffer_401),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_41),
	.datad(out_data_buffer_411),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_42),
	.datad(out_data_buffer_421),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_43),
	.datad(out_data_buffer_431),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_44),
	.datad(out_data_buffer_441),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_45),
	.datad(out_data_buffer_451),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_46),
	.datad(out_data_buffer_461),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[47] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_47),
	.datad(out_data_buffer_471),
	.cin(gnd),
	.combout(src_data_47),
	.cout());
defparam \src_data[47] .lut_mask = 16'hFFFE;
defparam \src_data[47] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_107),
	.datad(out_data_buffer_1071),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0] .lut_mask = 16'hFFFE;
defparam \src_payload[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(wire_pll7_clk_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(last_cycle),
	.datab(src_payload_0),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hACFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

endmodule

module usb_system_altera_merlin_arbitrator_3 (
	clk,
	reset,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	grant_0,
	update_grant,
	grant_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
output 	grant_0;
input 	update_grant;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~4_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~5_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(out_valid1),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(out_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~4 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(update_grant),
	.datad(out_valid),
	.cin(gnd),
	.combout(\top_priority_reg[0]~4_combout ),
	.cout());
defparam \top_priority_reg[0]~4 .lut_mask = 16'hFFF6;
defparam \top_priority_reg[0]~4 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~5 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~5_combout ),
	.cout());
defparam \top_priority_reg[0]~5 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~5 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module usb_system_usb_system_mm_interconnect_0_router (
	W_alu_result_7,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_12,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_8,
	W_alu_result_6,
	W_alu_result_24,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_3,
	Equal1,
	Equal3,
	Equal6,
	d_read,
	read_accepted,
	Equal2,
	always1,
	Equal11,
	uav_read,
	always11,
	Equal9,
	Equal91,
	always12,
	Equal5,
	Equal31,
	Equal7,
	Equal61,
	always13,
	Equal12,
	always14)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_12;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_8;
input 	W_alu_result_6;
input 	W_alu_result_24;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_28;
input 	W_alu_result_27;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_3;
output 	Equal1;
output 	Equal3;
output 	Equal6;
input 	d_read;
input 	read_accepted;
output 	Equal2;
output 	always1;
output 	Equal11;
input 	uav_read;
output 	always11;
output 	Equal9;
output 	Equal91;
output 	always12;
output 	Equal5;
output 	Equal31;
output 	Equal7;
output 	Equal61;
output 	always13;
output 	Equal12;
output 	always14;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal3~0_combout ;
wire \Equal3~1_combout ;
wire \Equal3~2_combout ;
wire \Equal2~2_combout ;
wire \Equal3~3_combout ;
wire \Equal1~1_combout ;
wire \Equal2~3_combout ;
wire \Equal2~4_combout ;
wire \Equal3~5_combout ;
wire \always1~7_combout ;
wire \Equal6~1_combout ;


cycloneive_lcell_comb \Equal1~0 (
	.dataa(W_alu_result_28),
	.datab(W_alu_result_27),
	.datac(W_alu_result_26),
	.datad(W_alu_result_25),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hBFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~4 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\Equal3~3_combout ),
	.cin(gnd),
	.combout(Equal3),
	.cout());
defparam \Equal3~4 .lut_mask = 16'hFFFE;
defparam \Equal3~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(W_alu_result_7),
	.datab(Equal3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~0 .lut_mask = 16'hEEEE;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~5 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Equal2~3_combout ),
	.datad(\Equal2~4_combout ),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~5 .lut_mask = 16'hFFFE;
defparam \Equal2~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~2 (
	.dataa(W_alu_result_5),
	.datab(d_read),
	.datac(W_alu_result_4),
	.datad(read_accepted),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~2 .lut_mask = 16'hEFFF;
defparam \always1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(W_alu_result_23),
	.datab(W_alu_result_22),
	.datac(W_alu_result_24),
	.datad(Equal1),
	.cin(gnd),
	.combout(Equal11),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hFEFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~3 (
	.dataa(W_alu_result_5),
	.datab(W_alu_result_3),
	.datac(uav_read),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(always11),
	.cout());
defparam \always1~3 .lut_mask = 16'hFEFF;
defparam \always1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal9~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_5),
	.datac(gnd),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(Equal9),
	.cout());
defparam \Equal9~0 .lut_mask = 16'hEEFF;
defparam \Equal9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal9~1 (
	.dataa(W_alu_result_7),
	.datab(Equal3),
	.datac(Equal9),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal91),
	.cout());
defparam \Equal9~1 .lut_mask = 16'hFEFE;
defparam \Equal9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~4 (
	.dataa(\Equal1~1_combout ),
	.datab(\Equal2~3_combout ),
	.datac(\Equal3~5_combout ),
	.datad(\always1~7_combout ),
	.cin(gnd),
	.combout(always12),
	.cout());
defparam \always1~4 .lut_mask = 16'hFFFE;
defparam \always1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_5),
	.datac(Equal3),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(Equal5),
	.cout());
defparam \Equal5~0 .lut_mask = 16'hFEFF;
defparam \Equal5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~6 (
	.dataa(W_alu_result_4),
	.datab(Equal3),
	.datac(W_alu_result_5),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(Equal31),
	.cout());
defparam \Equal3~6 .lut_mask = 16'hEFFF;
defparam \Equal3~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal7~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_7),
	.datac(Equal3),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(Equal7),
	.cout());
defparam \Equal7~0 .lut_mask = 16'hFEFF;
defparam \Equal7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~2 (
	.dataa(\Equal1~1_combout ),
	.datab(\Equal2~3_combout ),
	.datac(\Equal3~5_combout ),
	.datad(\Equal6~1_combout ),
	.cin(gnd),
	.combout(Equal61),
	.cout());
defparam \Equal6~2 .lut_mask = 16'hFFFE;
defparam \Equal6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~5 (
	.dataa(Equal3),
	.datab(always1),
	.datac(gnd),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(always13),
	.cout());
defparam \always1~5 .lut_mask = 16'hEEFF;
defparam \always1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_23),
	.datad(W_alu_result_22),
	.cin(gnd),
	.combout(Equal12),
	.cout());
defparam \Equal1~3 .lut_mask = 16'h0FFF;
defparam \Equal1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~6 (
	.dataa(W_alu_result_7),
	.datab(Equal3),
	.datac(always11),
	.datad(gnd),
	.cin(gnd),
	.combout(always14),
	.cout());
defparam \always1~6 .lut_mask = 16'hFEFE;
defparam \always1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_14),
	.datad(W_alu_result_13),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h0FFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_18),
	.datad(W_alu_result_17),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'h0FFF;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(W_alu_result_12),
	.datab(W_alu_result_11),
	.datac(W_alu_result_10),
	.datad(W_alu_result_9),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'hBFFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~1 (
	.dataa(W_alu_result_23),
	.datab(W_alu_result_22),
	.datac(W_alu_result_8),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
defparam \Equal3~1 .lut_mask = 16'h7FFF;
defparam \Equal3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~2 (
	.dataa(W_alu_result_16),
	.datab(W_alu_result_15),
	.datac(\Equal3~0_combout ),
	.datad(\Equal3~1_combout ),
	.cin(gnd),
	.combout(\Equal3~2_combout ),
	.cout());
defparam \Equal3~2 .lut_mask = 16'hFFF7;
defparam \Equal3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~2 (
	.dataa(W_alu_result_24),
	.datab(W_alu_result_21),
	.datac(W_alu_result_20),
	.datad(W_alu_result_19),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hBFFF;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~3 (
	.dataa(\Equal2~2_combout ),
	.datab(Equal1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal3~3_combout ),
	.cout());
defparam \Equal3~3 .lut_mask = 16'hEEEE;
defparam \Equal3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(Equal1),
	.datab(gnd),
	.datac(W_alu_result_23),
	.datad(W_alu_result_22),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hAFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~3 (
	.dataa(\Equal2~2_combout ),
	.datab(\Equal2~1_combout ),
	.datac(W_alu_result_16),
	.datad(W_alu_result_15),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
defparam \Equal2~3 .lut_mask = 16'hEFFF;
defparam \Equal2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~4 (
	.dataa(W_alu_result_11),
	.datab(gnd),
	.datac(gnd),
	.datad(W_alu_result_12),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
defparam \Equal2~4 .lut_mask = 16'hAAFF;
defparam \Equal2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~5 (
	.dataa(\Equal3~0_combout ),
	.datab(gnd),
	.datac(W_alu_result_8),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\Equal3~5_combout ),
	.cout());
defparam \Equal3~5 .lut_mask = 16'hAFFF;
defparam \Equal3~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~7 (
	.dataa(W_alu_result_14),
	.datab(W_alu_result_13),
	.datac(W_alu_result_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~7_combout ),
	.cout());
defparam \always1~7 .lut_mask = 16'h7F7F;
defparam \always1~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~1 (
	.dataa(W_alu_result_7),
	.datab(W_alu_result_4),
	.datac(W_alu_result_5),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\Equal6~1_combout ),
	.cout());
defparam \Equal6~1 .lut_mask = 16'hFFBF;
defparam \Equal6~1 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_router_001 (
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	Equal1,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_5,
	F_pc_6,
	F_pc_4,
	Equal2,
	F_pc_1,
	F_pc_3,
	i_read,
	read_accepted,
	F_pc_2,
	always1,
	Equal21,
	always11,
	Equal11)/* synthesis synthesis_greybox=1 */;
input 	F_pc_26;
input 	F_pc_25;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
output 	Equal1;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_5;
input 	F_pc_6;
input 	F_pc_4;
output 	Equal2;
input 	F_pc_1;
input 	F_pc_3;
input 	i_read;
input 	read_accepted;
input 	F_pc_2;
output 	always1;
output 	Equal21;
output 	always11;
output 	Equal11;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \Equal1~3_combout ;
wire \Equal2~0_combout ;
wire \always1~0_combout ;


cycloneive_lcell_comb \Equal1~4 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Equal1~2_combout ),
	.datad(\Equal1~3_combout ),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~4 .lut_mask = 16'hFFFE;
defparam \Equal1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(\Equal2~0_combout ),
	.datab(F_pc_5),
	.datac(F_pc_6),
	.datad(F_pc_4),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hEFFF;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~1 (
	.dataa(F_pc_1),
	.datab(\always1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~1 .lut_mask = 16'hEEEE;
defparam \always1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~2 (
	.dataa(Equal1),
	.datab(Equal2),
	.datac(F_pc_2),
	.datad(F_pc_3),
	.cin(gnd),
	.combout(Equal21),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hFEFF;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~2 (
	.dataa(Equal1),
	.datab(Equal2),
	.datac(F_pc_1),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(always11),
	.cout());
defparam \always1~2 .lut_mask = 16'hFFFE;
defparam \always1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~5 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(Equal1),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(Equal11),
	.cout());
defparam \Equal1~5 .lut_mask = 16'hAFFF;
defparam \Equal1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(F_pc_26),
	.datab(F_pc_25),
	.datac(F_pc_24),
	.datad(F_pc_23),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(F_pc_22),
	.datab(F_pc_21),
	.datac(F_pc_20),
	.datad(F_pc_19),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hBFFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(F_pc_18),
	.datab(F_pc_17),
	.datac(F_pc_16),
	.datad(F_pc_15),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'h7FFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~3 (
	.dataa(F_pc_14),
	.datab(F_pc_13),
	.datac(F_pc_12),
	.datad(F_pc_11),
	.cin(gnd),
	.combout(\Equal1~3_combout ),
	.cout());
defparam \Equal1~3 .lut_mask = 16'h7FFF;
defparam \Equal1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(F_pc_10),
	.datab(F_pc_9),
	.datac(F_pc_8),
	.datad(F_pc_7),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hBFFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(F_pc_3),
	.datab(i_read),
	.datac(read_accepted),
	.datad(F_pc_2),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hBFFF;
defparam \always1~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_router_003_3 (
	mem_86_0,
	mem_68_0,
	always0)/* synthesis synthesis_greybox=1 */;
input 	mem_86_0;
input 	mem_68_0;
output 	always0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \always0~0 (
	.dataa(mem_86_0),
	.datab(mem_68_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hEEEE;
defparam \always0~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_rsp_demux_001 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_rsp_demux_001_1 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_rsp_demux_001_2 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_rsp_demux_001_3 (
	mem_86_0,
	mem_68_0,
	in_data_toggle,
	dreg_0,
	in_data_toggle1,
	dreg_01,
	always0,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	mem_86_0;
input 	mem_68_0;
input 	in_data_toggle;
input 	dreg_0;
input 	in_data_toggle1;
input 	dreg_01;
input 	always0;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;


cycloneive_lcell_comb \WideOr0~1 (
	.dataa(\WideOr0~0_combout ),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(always0),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hBEFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(mem_86_0),
	.datab(mem_68_0),
	.datac(in_data_toggle),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_rsp_mux (
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	out_valid,
	read_latency_shift_reg_02,
	mem_86_0,
	mem_68_0,
	src0_valid,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	mem_86_01,
	mem_68_01,
	src0_valid1,
	read_latency_shift_reg_05,
	mem_86_02,
	mem_68_02,
	read_latency_shift_reg_06,
	read_latency_shift_reg_07,
	out_data_toggle_flopped,
	dreg_0,
	WideOr11,
	src0_valid2,
	out_valid1,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_1,
	av_readdata_pre_11,
	av_readdata_pre_2,
	av_readdata_pre_30,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_02,
	out_payload_0,
	av_readdata_pre_03,
	av_readdata_pre_04,
	av_readdata_pre_05,
	av_readdata_pre_06,
	out_data_buffer_0,
	src_data_0,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_111,
	av_readdata_pre_13,
	av_readdata_pre_161,
	av_readdata_pre_12,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_201,
	av_readdata_pre_181,
	av_readdata_pre_191,
	av_readdata_pre_171,
	av_readdata_pre_211,
	av_readdata_pre_110,
	out_payload_1,
	av_readdata_pre_112,
	av_readdata_pre_113,
	av_readdata_pre_114,
	av_readdata_pre_115,
	out_data_buffer_1,
	src_data_1,
	src_payload,
	av_readdata_pre_24,
	out_payload_2,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_data_2,
	av_readdata_pre_27,
	av_readdata_pre_28,
	out_data_buffer_2,
	av_readdata_pre_31,
	av_readdata_pre_32,
	src_data_3,
	av_readdata_pre_33,
	out_payload_3,
	av_readdata_pre_34,
	av_readdata_pre_35,
	out_data_buffer_3,
	src_data_31,
	av_readdata_pre_41,
	out_payload_4,
	av_readdata_pre_42,
	av_readdata_pre_43,
	src_data_4,
	av_readdata_pre_44,
	av_readdata_pre_45,
	out_data_buffer_4,
	av_readdata_pre_51,
	out_payload_5,
	av_readdata_pre_52,
	av_readdata_pre_53,
	src_data_5,
	av_readdata_pre_54,
	av_readdata_pre_55,
	out_data_buffer_5,
	av_readdata_pre_61,
	out_payload_6,
	av_readdata_pre_62,
	av_readdata_pre_63,
	src_data_6,
	av_readdata_pre_64,
	av_readdata_pre_65,
	out_data_buffer_6,
	av_readdata_pre_71,
	out_payload_7,
	av_readdata_pre_72,
	av_readdata_pre_73,
	src_data_7,
	av_readdata_pre_74,
	av_readdata_pre_75,
	out_data_buffer_7,
	av_readdata_pre_81,
	av_readdata_pre_82,
	out_data_buffer_8,
	av_readdata_pre_83,
	out_payload_8,
	src_data_8,
	av_readdata_pre_91,
	av_readdata_pre_92,
	av_readdata_pre_93,
	out_payload_9,
	out_data_buffer_9,
	src_data_9,
	av_readdata_pre_101,
	out_payload_10,
	av_readdata_pre_102,
	av_readdata_pre_103,
	out_data_buffer_10,
	src_data_10,
	av_readdata_pre_116,
	out_payload_11,
	out_data_buffer_11,
	av_readdata_pre_117,
	src_data_11,
	av_readdata_pre_121,
	out_payload_12,
	av_readdata_pre_122,
	av_readdata_pre_123,
	out_data_buffer_12,
	src_data_12,
	av_readdata_pre_131,
	av_readdata_pre_132,
	av_readdata_pre_133,
	out_payload_13,
	out_data_buffer_13,
	src_data_13,
	av_readdata_pre_141,
	out_payload_14,
	av_readdata_pre_142,
	av_readdata_pre_143,
	out_data_buffer_14,
	src_data_14,
	av_readdata_pre_151,
	av_readdata_pre_152,
	out_data_buffer_15,
	av_readdata_pre_153,
	out_payload_15,
	src_data_15,
	av_readdata_pre_162,
	out_data_buffer_16,
	av_readdata_pre_163,
	src_data_16,
	av_readdata_pre_172,
	out_data_buffer_17,
	av_readdata_pre_173,
	src_data_17,
	out_data_buffer_18,
	src_payload1,
	out_data_buffer_23,
	src_payload2,
	out_data_buffer_22,
	src_payload3,
	out_data_buffer_21,
	src_payload4,
	out_data_buffer_20,
	src_payload5,
	out_data_buffer_19,
	src_payload6,
	src_data_21,
	src_data_41,
	src_data_51,
	src_data_61,
	src_data_71)/* synthesis synthesis_greybox=1 */;
input 	av_readdata_pre_16;
input 	av_readdata_pre_17;
input 	av_readdata_pre_18;
input 	av_readdata_pre_22;
input 	av_readdata_pre_21;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	out_valid;
input 	read_latency_shift_reg_02;
input 	mem_86_0;
input 	mem_68_0;
input 	src0_valid;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
input 	mem_86_01;
input 	mem_68_01;
input 	src0_valid1;
input 	read_latency_shift_reg_05;
input 	mem_86_02;
input 	mem_68_02;
input 	read_latency_shift_reg_06;
input 	read_latency_shift_reg_07;
input 	out_data_toggle_flopped;
input 	dreg_0;
output 	WideOr11;
input 	src0_valid2;
input 	out_valid1;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	av_readdata_pre_2;
input 	av_readdata_pre_30;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_02;
input 	out_payload_0;
input 	av_readdata_pre_03;
input 	av_readdata_pre_04;
input 	av_readdata_pre_05;
input 	av_readdata_pre_06;
input 	out_data_buffer_0;
output 	src_data_0;
input 	av_readdata_pre_221;
input 	av_readdata_pre_23;
input 	av_readdata_pre_111;
input 	av_readdata_pre_13;
input 	av_readdata_pre_161;
input 	av_readdata_pre_12;
input 	av_readdata_pre_5;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_10;
input 	av_readdata_pre_9;
input 	av_readdata_pre_8;
input 	av_readdata_pre_7;
input 	av_readdata_pre_6;
input 	av_readdata_pre_201;
input 	av_readdata_pre_181;
input 	av_readdata_pre_191;
input 	av_readdata_pre_171;
input 	av_readdata_pre_211;
input 	av_readdata_pre_110;
input 	out_payload_1;
input 	av_readdata_pre_112;
input 	av_readdata_pre_113;
input 	av_readdata_pre_114;
input 	av_readdata_pre_115;
input 	out_data_buffer_1;
output 	src_data_1;
output 	src_payload;
input 	av_readdata_pre_24;
input 	out_payload_2;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
output 	src_data_2;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	out_data_buffer_2;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
output 	src_data_3;
input 	av_readdata_pre_33;
input 	out_payload_3;
input 	av_readdata_pre_34;
input 	av_readdata_pre_35;
input 	out_data_buffer_3;
output 	src_data_31;
input 	av_readdata_pre_41;
input 	out_payload_4;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
output 	src_data_4;
input 	av_readdata_pre_44;
input 	av_readdata_pre_45;
input 	out_data_buffer_4;
input 	av_readdata_pre_51;
input 	out_payload_5;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
output 	src_data_5;
input 	av_readdata_pre_54;
input 	av_readdata_pre_55;
input 	out_data_buffer_5;
input 	av_readdata_pre_61;
input 	out_payload_6;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
output 	src_data_6;
input 	av_readdata_pre_64;
input 	av_readdata_pre_65;
input 	out_data_buffer_6;
input 	av_readdata_pre_71;
input 	out_payload_7;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
output 	src_data_7;
input 	av_readdata_pre_74;
input 	av_readdata_pre_75;
input 	out_data_buffer_7;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
input 	out_data_buffer_8;
input 	av_readdata_pre_83;
input 	out_payload_8;
output 	src_data_8;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
input 	av_readdata_pre_93;
input 	out_payload_9;
input 	out_data_buffer_9;
output 	src_data_9;
input 	av_readdata_pre_101;
input 	out_payload_10;
input 	av_readdata_pre_102;
input 	av_readdata_pre_103;
input 	out_data_buffer_10;
output 	src_data_10;
input 	av_readdata_pre_116;
input 	out_payload_11;
input 	out_data_buffer_11;
input 	av_readdata_pre_117;
output 	src_data_11;
input 	av_readdata_pre_121;
input 	out_payload_12;
input 	av_readdata_pre_122;
input 	av_readdata_pre_123;
input 	out_data_buffer_12;
output 	src_data_12;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
input 	av_readdata_pre_133;
input 	out_payload_13;
input 	out_data_buffer_13;
output 	src_data_13;
input 	av_readdata_pre_141;
input 	out_payload_14;
input 	av_readdata_pre_142;
input 	av_readdata_pre_143;
input 	out_data_buffer_14;
output 	src_data_14;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
input 	out_data_buffer_15;
input 	av_readdata_pre_153;
input 	out_payload_15;
output 	src_data_15;
input 	av_readdata_pre_162;
input 	out_data_buffer_16;
input 	av_readdata_pre_163;
output 	src_data_16;
input 	av_readdata_pre_172;
input 	out_data_buffer_17;
input 	av_readdata_pre_173;
output 	src_data_17;
input 	out_data_buffer_18;
output 	src_payload1;
input 	out_data_buffer_23;
output 	src_payload2;
input 	out_data_buffer_22;
output 	src_payload3;
input 	out_data_buffer_21;
output 	src_payload4;
input 	out_data_buffer_20;
output 	src_payload5;
input 	out_data_buffer_19;
output 	src_payload6;
output 	src_data_21;
output 	src_data_41;
output 	src_data_51;
output 	src_data_61;
output 	src_data_71;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;
wire \WideOr1~2_combout ;
wire \src_data[0]~18_combout ;
wire \src_data[0]~19_combout ;
wire \src_data[0]~20_combout ;
wire \src_data[0]~21_combout ;
wire \src_data[0]~82_combout ;
wire \src_data[1]~22_combout ;
wire \src_data[1]~23_combout ;
wire \src_data[1]~24_combout ;
wire \src_data[1]~25_combout ;
wire \src_data[1]~83_combout ;
wire \src_payload~1_combout ;
wire \src_data[2]~26_combout ;
wire \src_data[2]~27_combout ;
wire \src_data[3]~31_combout ;
wire \src_data[3]~32_combout ;
wire \src_data[3]~33_combout ;
wire \src_payload~2_combout ;
wire \src_data[4]~35_combout ;
wire \src_data[4]~36_combout ;
wire \src_payload~3_combout ;
wire \src_data[5]~39_combout ;
wire \src_data[5]~40_combout ;
wire \src_payload~4_combout ;
wire \src_data[6]~43_combout ;
wire \src_data[6]~44_combout ;
wire \src_payload~5_combout ;
wire \src_data[7]~47_combout ;
wire \src_data[7]~48_combout ;
wire \src_data[8]~51_combout ;
wire \src_data[8]~52_combout ;
wire \src_payload~6_combout ;
wire \src_data[8]~53_combout ;
wire \src_data[9]~54_combout ;
wire \src_payload~7_combout ;
wire \src_data[9]~55_combout ;
wire \src_data[9]~89_combout ;
wire \src_data[10]~56_combout ;
wire \src_data[10]~57_combout ;
wire \src_data[10]~58_combout ;
wire \src_data[11]~60_combout ;
wire \src_data[11]~61_combout ;
wire \src_data[11]~62_combout ;
wire \src_data[12]~63_combout ;
wire \src_data[12]~64_combout ;
wire \src_data[12]~65_combout ;
wire \src_data[13]~67_combout ;
wire \src_payload~8_combout ;
wire \src_data[13]~68_combout ;
wire \src_data[13]~90_combout ;
wire \src_data[14]~69_combout ;
wire \src_data[14]~70_combout ;
wire \src_data[14]~71_combout ;
wire \src_data[15]~73_combout ;
wire \src_data[15]~74_combout ;
wire \src_payload~9_combout ;
wire \src_data[15]~75_combout ;
wire \src_data[16]~76_combout ;
wire \src_data[16]~77_combout ;
wire \src_data[17]~79_combout ;
wire \src_data[17]~80_combout ;
wire \src_data[17]~81_combout ;
wire \src_payload~10_combout ;
wire \src_payload~13_combout ;
wire \src_payload~15_combout ;
wire \src_payload~17_combout ;
wire \src_payload~19_combout ;
wire \src_data[2]~29_combout ;
wire \src_data[4]~38_combout ;
wire \src_data[5]~42_combout ;
wire \src_data[6]~46_combout ;
wire \src_data[7]~50_combout ;


cycloneive_lcell_comb WideOr1(
	.dataa(read_latency_shift_reg_01),
	.datab(\WideOr1~0_combout ),
	.datac(\WideOr1~1_combout ),
	.datad(\WideOr1~2_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0] (
	.dataa(\src_data[0]~18_combout ),
	.datab(\src_data[0]~19_combout ),
	.datac(\src_data[0]~20_combout ),
	.datad(\src_data[0]~82_combout ),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0] .lut_mask = 16'hFFFE;
defparam \src_data[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1] (
	.dataa(\src_data[1]~22_combout ),
	.datab(\src_data[1]~23_combout ),
	.datac(\src_data[1]~24_combout ),
	.datad(\src_data[1]~83_combout ),
	.cin(gnd),
	.combout(src_data_1),
	.cout());
defparam \src_data[1] .lut_mask = 16'hFFFE;
defparam \src_data[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_02),
	.datab(av_readdata_pre_30),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEFFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~28 (
	.dataa(src_payload),
	.datab(\src_payload~1_combout ),
	.datac(\src_data[2]~26_combout ),
	.datad(\src_data[2]~27_combout ),
	.cin(gnd),
	.combout(src_data_2),
	.cout());
defparam \src_data[2]~28 .lut_mask = 16'hFFFE;
defparam \src_data[2]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~30 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_31),
	.datad(av_readdata_pre_32),
	.cin(gnd),
	.combout(src_data_3),
	.cout());
defparam \src_data[3]~30 .lut_mask = 16'hFFFE;
defparam \src_data[3]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~34 (
	.dataa(\src_data[3]~32_combout ),
	.datab(\src_data[3]~33_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_3),
	.cin(gnd),
	.combout(src_data_31),
	.cout());
defparam \src_data[3]~34 .lut_mask = 16'hFFFE;
defparam \src_data[3]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~37 (
	.dataa(src_payload),
	.datab(\src_payload~2_combout ),
	.datac(\src_data[4]~35_combout ),
	.datad(\src_data[4]~36_combout ),
	.cin(gnd),
	.combout(src_data_4),
	.cout());
defparam \src_data[4]~37 .lut_mask = 16'hFFFE;
defparam \src_data[4]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~41 (
	.dataa(src_payload),
	.datab(\src_payload~3_combout ),
	.datac(\src_data[5]~39_combout ),
	.datad(\src_data[5]~40_combout ),
	.cin(gnd),
	.combout(src_data_5),
	.cout());
defparam \src_data[5]~41 .lut_mask = 16'hFFFE;
defparam \src_data[5]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~45 (
	.dataa(src_payload),
	.datab(\src_payload~4_combout ),
	.datac(\src_data[6]~43_combout ),
	.datad(\src_data[6]~44_combout ),
	.cin(gnd),
	.combout(src_data_6),
	.cout());
defparam \src_data[6]~45 .lut_mask = 16'hFFFE;
defparam \src_data[6]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~49 (
	.dataa(src_payload),
	.datab(\src_payload~5_combout ),
	.datac(\src_data[7]~47_combout ),
	.datad(\src_data[7]~48_combout ),
	.cin(gnd),
	.combout(src_data_7),
	.cout());
defparam \src_data[7]~49 .lut_mask = 16'hFFFE;
defparam \src_data[7]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8] (
	.dataa(\src_data[8]~51_combout ),
	.datab(\src_data[8]~52_combout ),
	.datac(\src_payload~6_combout ),
	.datad(\src_data[8]~53_combout ),
	.cin(gnd),
	.combout(src_data_8),
	.cout());
defparam \src_data[8] .lut_mask = 16'hFFFE;
defparam \src_data[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9] (
	.dataa(src_payload),
	.datab(\src_data[9]~54_combout ),
	.datac(\src_payload~7_combout ),
	.datad(\src_data[9]~89_combout ),
	.cin(gnd),
	.combout(src_data_9),
	.cout());
defparam \src_data[9] .lut_mask = 16'hFFFE;
defparam \src_data[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~59 (
	.dataa(\src_data[10]~57_combout ),
	.datab(\src_data[10]~58_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_10),
	.cin(gnd),
	.combout(src_data_10),
	.cout());
defparam \src_data[10]~59 .lut_mask = 16'hFFFE;
defparam \src_data[10]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11] (
	.dataa(\src_data[11]~62_combout ),
	.datab(read_latency_shift_reg_01),
	.datac(av_readdata_pre_117),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_11),
	.cout());
defparam \src_data[11] .lut_mask = 16'hFEFE;
defparam \src_data[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~66 (
	.dataa(\src_data[12]~64_combout ),
	.datab(\src_data[12]~65_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_12),
	.cin(gnd),
	.combout(src_data_12),
	.cout());
defparam \src_data[12]~66 .lut_mask = 16'hFFFE;
defparam \src_data[12]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13] (
	.dataa(src_payload),
	.datab(\src_data[13]~67_combout ),
	.datac(\src_payload~8_combout ),
	.datad(\src_data[13]~90_combout ),
	.cin(gnd),
	.combout(src_data_13),
	.cout());
defparam \src_data[13] .lut_mask = 16'hFFFE;
defparam \src_data[13] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~72 (
	.dataa(\src_data[14]~70_combout ),
	.datab(\src_data[14]~71_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_14),
	.cin(gnd),
	.combout(src_data_14),
	.cout());
defparam \src_data[14]~72 .lut_mask = 16'hFFFE;
defparam \src_data[14]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15] (
	.dataa(\src_data[15]~73_combout ),
	.datab(\src_data[15]~74_combout ),
	.datac(\src_payload~9_combout ),
	.datad(\src_data[15]~75_combout ),
	.cin(gnd),
	.combout(src_data_15),
	.cout());
defparam \src_data[15] .lut_mask = 16'hFFFE;
defparam \src_data[15] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~78 (
	.dataa(\src_data[16]~76_combout ),
	.datab(\src_data[16]~77_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_161),
	.cin(gnd),
	.combout(src_data_16),
	.cout());
defparam \src_data[16]~78 .lut_mask = 16'hFFFE;
defparam \src_data[16]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17] (
	.dataa(\src_data[17]~81_combout ),
	.datab(read_latency_shift_reg_01),
	.datac(av_readdata_pre_173),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_17),
	.cout());
defparam \src_data[17] .lut_mask = 16'hFEFE;
defparam \src_data[17] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(\src_payload~10_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_181),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hFEFE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(src0_valid1),
	.datab(out_valid1),
	.datac(out_data_buffer_23),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hFFFE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(src_payload),
	.datab(\src_payload~13_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_221),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hFFFE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(\src_payload~15_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_211),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hFEFE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(\src_payload~17_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_201),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hFEFE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(src_payload),
	.datab(\src_payload~19_combout ),
	.datac(src0_valid1),
	.datad(av_readdata_pre_191),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hFFFE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~84 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[2]~29_combout ),
	.datad(out_data_buffer_2),
	.cin(gnd),
	.combout(src_data_21),
	.cout());
defparam \src_data[2]~84 .lut_mask = 16'hFFF6;
defparam \src_data[2]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~85 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[4]~38_combout ),
	.datad(out_data_buffer_4),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[4]~85 .lut_mask = 16'hFFF6;
defparam \src_data[4]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~86 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[5]~42_combout ),
	.datad(out_data_buffer_5),
	.cin(gnd),
	.combout(src_data_51),
	.cout());
defparam \src_data[5]~86 .lut_mask = 16'hFFF6;
defparam \src_data[5]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~87 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[6]~46_combout ),
	.datad(out_data_buffer_6),
	.cin(gnd),
	.combout(src_data_61),
	.cout());
defparam \src_data[6]~87 .lut_mask = 16'hFFF6;
defparam \src_data[6]~87 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~88 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[7]~50_combout ),
	.datad(out_data_buffer_7),
	.cin(gnd),
	.combout(src_data_71),
	.cout());
defparam \src_data[7]~88 .lut_mask = 16'hFFF6;
defparam \src_data[7]~88 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(out_valid),
	.datab(src0_valid),
	.datac(read_latency_shift_reg_03),
	.datad(src0_valid1),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~1 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_05),
	.datac(mem_86_02),
	.datad(mem_68_02),
	.cin(gnd),
	.combout(\WideOr1~1_combout ),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'hEFFF;
defparam \WideOr1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~2 (
	.dataa(read_latency_shift_reg_06),
	.datab(read_latency_shift_reg_07),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\WideOr1~2_combout ),
	.cout());
defparam \WideOr1~2 .lut_mask = 16'hEFFE;
defparam \WideOr1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~18 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(av_readdata_pre_0),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(\src_data[0]~18_combout ),
	.cout());
defparam \src_data[0]~18 .lut_mask = 16'hFFFE;
defparam \src_data[0]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~19 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_02),
	.datad(out_payload_0),
	.cin(gnd),
	.combout(\src_data[0]~19_combout ),
	.cout());
defparam \src_data[0]~19 .lut_mask = 16'hFFFE;
defparam \src_data[0]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~20 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_03),
	.datad(av_readdata_pre_04),
	.cin(gnd),
	.combout(\src_data[0]~20_combout ),
	.cout());
defparam \src_data[0]~20 .lut_mask = 16'hFFFE;
defparam \src_data[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~21 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_05),
	.datad(av_readdata_pre_06),
	.cin(gnd),
	.combout(\src_data[0]~21_combout ),
	.cout());
defparam \src_data[0]~21 .lut_mask = 16'hFFFE;
defparam \src_data[0]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~82 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[0]~21_combout ),
	.datad(out_data_buffer_0),
	.cin(gnd),
	.combout(\src_data[0]~82_combout ),
	.cout());
defparam \src_data[0]~82 .lut_mask = 16'hFFF6;
defparam \src_data[0]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~22 (
	.dataa(src0_valid1),
	.datab(src0_valid2),
	.datac(av_readdata_pre_1),
	.datad(av_readdata_pre_11),
	.cin(gnd),
	.combout(\src_data[1]~22_combout ),
	.cout());
defparam \src_data[1]~22 .lut_mask = 16'hFFFE;
defparam \src_data[1]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~23 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_110),
	.datad(out_payload_1),
	.cin(gnd),
	.combout(\src_data[1]~23_combout ),
	.cout());
defparam \src_data[1]~23 .lut_mask = 16'hFFFE;
defparam \src_data[1]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~24 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_112),
	.datad(av_readdata_pre_113),
	.cin(gnd),
	.combout(\src_data[1]~24_combout ),
	.cout());
defparam \src_data[1]~24 .lut_mask = 16'hFFFE;
defparam \src_data[1]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~25 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_114),
	.datad(av_readdata_pre_115),
	.cin(gnd),
	.combout(\src_data[1]~25_combout ),
	.cout());
defparam \src_data[1]~25 .lut_mask = 16'hFFFE;
defparam \src_data[1]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~83 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[1]~25_combout ),
	.datad(out_data_buffer_1),
	.cin(gnd),
	.combout(\src_data[1]~83_combout ),
	.cout());
defparam \src_data[1]~83 .lut_mask = 16'hFFF6;
defparam \src_data[1]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_2),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~1_combout ),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEFFF;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~26 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_24),
	.datad(out_payload_2),
	.cin(gnd),
	.combout(\src_data[2]~26_combout ),
	.cout());
defparam \src_data[2]~26 .lut_mask = 16'hFFFE;
defparam \src_data[2]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~27 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_25),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\src_data[2]~27_combout ),
	.cout());
defparam \src_data[2]~27 .lut_mask = 16'hFFFE;
defparam \src_data[2]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~31 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_33),
	.datad(out_payload_3),
	.cin(gnd),
	.combout(\src_data[3]~31_combout ),
	.cout());
defparam \src_data[3]~31 .lut_mask = 16'hFFFE;
defparam \src_data[3]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~32 (
	.dataa(\src_data[3]~31_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[3]~32_combout ),
	.cout());
defparam \src_data[3]~32 .lut_mask = 16'hFEFE;
defparam \src_data[3]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~33 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_34),
	.datad(av_readdata_pre_35),
	.cin(gnd),
	.combout(\src_data[3]~33_combout ),
	.cout());
defparam \src_data[3]~33 .lut_mask = 16'hFFFE;
defparam \src_data[3]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_4),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~2_combout ),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEFFF;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~35 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_41),
	.datad(out_payload_4),
	.cin(gnd),
	.combout(\src_data[4]~35_combout ),
	.cout());
defparam \src_data[4]~35 .lut_mask = 16'hFFFE;
defparam \src_data[4]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~36 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_42),
	.datad(av_readdata_pre_43),
	.cin(gnd),
	.combout(\src_data[4]~36_combout ),
	.cout());
defparam \src_data[4]~36 .lut_mask = 16'hFFFE;
defparam \src_data[4]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_5),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~3_combout ),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEFFF;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~39 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_51),
	.datad(out_payload_5),
	.cin(gnd),
	.combout(\src_data[5]~39_combout ),
	.cout());
defparam \src_data[5]~39 .lut_mask = 16'hFFFE;
defparam \src_data[5]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~40 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_52),
	.datad(av_readdata_pre_53),
	.cin(gnd),
	.combout(\src_data[5]~40_combout ),
	.cout());
defparam \src_data[5]~40 .lut_mask = 16'hFFFE;
defparam \src_data[5]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_6),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~4_combout ),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEFFF;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~43 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_61),
	.datad(out_payload_6),
	.cin(gnd),
	.combout(\src_data[6]~43_combout ),
	.cout());
defparam \src_data[6]~43 .lut_mask = 16'hFFFE;
defparam \src_data[6]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~44 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_62),
	.datad(av_readdata_pre_63),
	.cin(gnd),
	.combout(\src_data[6]~44_combout ),
	.cout());
defparam \src_data[6]~44 .lut_mask = 16'hFFFE;
defparam \src_data[6]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_7),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~5_combout ),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEFFF;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~47 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_71),
	.datad(out_payload_7),
	.cin(gnd),
	.combout(\src_data[7]~47_combout ),
	.cout());
defparam \src_data[7]~47 .lut_mask = 16'hFFFE;
defparam \src_data[7]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~48 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_06),
	.datac(av_readdata_pre_72),
	.datad(av_readdata_pre_73),
	.cin(gnd),
	.combout(\src_data[7]~48_combout ),
	.cout());
defparam \src_data[7]~48 .lut_mask = 16'hFFFE;
defparam \src_data[7]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~51 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_81),
	.datad(av_readdata_pre_82),
	.cin(gnd),
	.combout(\src_data[8]~51_combout ),
	.cout());
defparam \src_data[8]~51 .lut_mask = 16'hFFFE;
defparam \src_data[8]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~52 (
	.dataa(src_payload),
	.datab(src0_valid1),
	.datac(av_readdata_pre_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[8]~52_combout ),
	.cout());
defparam \src_data[8]~52 .lut_mask = 16'hFEFE;
defparam \src_data[8]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(out_data_buffer_8),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\src_payload~6_combout ),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hAFFA;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~53 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_83),
	.datad(out_payload_8),
	.cin(gnd),
	.combout(\src_data[8]~53_combout ),
	.cout());
defparam \src_data[8]~53 .lut_mask = 16'hFFFE;
defparam \src_data[8]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~54 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_91),
	.datad(av_readdata_pre_92),
	.cin(gnd),
	.combout(\src_data[9]~54_combout ),
	.cout());
defparam \src_data[9]~54 .lut_mask = 16'hFFFE;
defparam \src_data[9]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_9),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~7_combout ),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEFFF;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~55 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_93),
	.datad(out_payload_9),
	.cin(gnd),
	.combout(\src_data[9]~55_combout ),
	.cout());
defparam \src_data[9]~55 .lut_mask = 16'hFFFE;
defparam \src_data[9]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~89 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[9]~55_combout ),
	.datad(out_data_buffer_9),
	.cin(gnd),
	.combout(\src_data[9]~89_combout ),
	.cout());
defparam \src_data[9]~89 .lut_mask = 16'hFFF6;
defparam \src_data[9]~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~56 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_101),
	.datad(out_payload_10),
	.cin(gnd),
	.combout(\src_data[10]~56_combout ),
	.cout());
defparam \src_data[10]~56 .lut_mask = 16'hFFFE;
defparam \src_data[10]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~57 (
	.dataa(\src_data[10]~56_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[10]~57_combout ),
	.cout());
defparam \src_data[10]~57 .lut_mask = 16'hFEFE;
defparam \src_data[10]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~58 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_102),
	.datad(av_readdata_pre_103),
	.cin(gnd),
	.combout(\src_data[10]~58_combout ),
	.cout());
defparam \src_data[10]~58 .lut_mask = 16'hFFFE;
defparam \src_data[10]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~60 (
	.dataa(src_payload),
	.datab(src0_valid1),
	.datac(av_readdata_pre_111),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[11]~60_combout ),
	.cout());
defparam \src_data[11]~60 .lut_mask = 16'hFEFE;
defparam \src_data[11]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~61 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_116),
	.datad(out_payload_11),
	.cin(gnd),
	.combout(\src_data[11]~61_combout ),
	.cout());
defparam \src_data[11]~61 .lut_mask = 16'hFFFE;
defparam \src_data[11]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~62 (
	.dataa(\src_data[11]~60_combout ),
	.datab(\src_data[11]~61_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_11),
	.cin(gnd),
	.combout(\src_data[11]~62_combout ),
	.cout());
defparam \src_data[11]~62 .lut_mask = 16'hFFFE;
defparam \src_data[11]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~63 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_121),
	.datad(out_payload_12),
	.cin(gnd),
	.combout(\src_data[12]~63_combout ),
	.cout());
defparam \src_data[12]~63 .lut_mask = 16'hFFFE;
defparam \src_data[12]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~64 (
	.dataa(\src_data[12]~63_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[12]~64_combout ),
	.cout());
defparam \src_data[12]~64 .lut_mask = 16'hFEFE;
defparam \src_data[12]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~65 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_122),
	.datad(av_readdata_pre_123),
	.cin(gnd),
	.combout(\src_data[12]~65_combout ),
	.cout());
defparam \src_data[12]~65 .lut_mask = 16'hFFFE;
defparam \src_data[12]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~67 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_131),
	.datad(av_readdata_pre_132),
	.cin(gnd),
	.combout(\src_data[13]~67_combout ),
	.cout());
defparam \src_data[13]~67 .lut_mask = 16'hFFFE;
defparam \src_data[13]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_13),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(\src_payload~8_combout ),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEFFF;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~68 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_133),
	.datad(out_payload_13),
	.cin(gnd),
	.combout(\src_data[13]~68_combout ),
	.cout());
defparam \src_data[13]~68 .lut_mask = 16'hFFFE;
defparam \src_data[13]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~90 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[13]~68_combout ),
	.datad(out_data_buffer_13),
	.cin(gnd),
	.combout(\src_data[13]~90_combout ),
	.cout());
defparam \src_data[13]~90 .lut_mask = 16'hFFF6;
defparam \src_data[13]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~69 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_141),
	.datad(out_payload_14),
	.cin(gnd),
	.combout(\src_data[14]~69_combout ),
	.cout());
defparam \src_data[14]~69 .lut_mask = 16'hFFFE;
defparam \src_data[14]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~70 (
	.dataa(\src_data[14]~69_combout ),
	.datab(src0_valid1),
	.datac(av_readdata_pre_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[14]~70_combout ),
	.cout());
defparam \src_data[14]~70 .lut_mask = 16'hFEFE;
defparam \src_data[14]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~71 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_142),
	.datad(av_readdata_pre_143),
	.cin(gnd),
	.combout(\src_data[14]~71_combout ),
	.cout());
defparam \src_data[14]~71 .lut_mask = 16'hFFFE;
defparam \src_data[14]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~73 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_151),
	.datad(av_readdata_pre_152),
	.cin(gnd),
	.combout(\src_data[15]~73_combout ),
	.cout());
defparam \src_data[15]~73 .lut_mask = 16'hFFFE;
defparam \src_data[15]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~74 (
	.dataa(src_payload),
	.datab(src0_valid1),
	.datac(av_readdata_pre_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[15]~74_combout ),
	.cout());
defparam \src_data[15]~74 .lut_mask = 16'hFEFE;
defparam \src_data[15]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(out_data_buffer_15),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\src_payload~9_combout ),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hAFFA;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~75 (
	.dataa(out_valid),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_153),
	.datad(out_payload_15),
	.cin(gnd),
	.combout(\src_data[15]~75_combout ),
	.cout());
defparam \src_data[15]~75 .lut_mask = 16'hFFFE;
defparam \src_data[15]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~76 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_162),
	.datad(av_readdata_pre_16),
	.cin(gnd),
	.combout(\src_data[16]~76_combout ),
	.cout());
defparam \src_data[16]~76 .lut_mask = 16'hFFFE;
defparam \src_data[16]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~77 (
	.dataa(read_latency_shift_reg_01),
	.datab(out_valid1),
	.datac(out_data_buffer_16),
	.datad(av_readdata_pre_163),
	.cin(gnd),
	.combout(\src_data[16]~77_combout ),
	.cout());
defparam \src_data[16]~77 .lut_mask = 16'hFFFE;
defparam \src_data[16]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~79 (
	.dataa(src_payload),
	.datab(src0_valid1),
	.datac(av_readdata_pre_171),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[17]~79_combout ),
	.cout());
defparam \src_data[17]~79 .lut_mask = 16'hFEFE;
defparam \src_data[17]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~80 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_172),
	.datad(av_readdata_pre_17),
	.cin(gnd),
	.combout(\src_data[17]~80_combout ),
	.cout());
defparam \src_data[17]~80 .lut_mask = 16'hFFFE;
defparam \src_data[17]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~81 (
	.dataa(\src_data[17]~79_combout ),
	.datab(\src_data[17]~80_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_17),
	.cin(gnd),
	.combout(\src_data[17]~81_combout ),
	.cout());
defparam \src_data[17]~81 .lut_mask = 16'hFFFE;
defparam \src_data[17]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(read_latency_shift_reg_03),
	.datab(out_valid1),
	.datac(out_data_buffer_18),
	.datad(av_readdata_pre_18),
	.cin(gnd),
	.combout(\src_payload~10_combout ),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hFFFE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(read_latency_shift_reg_03),
	.datab(out_valid1),
	.datac(out_data_buffer_22),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\src_payload~13_combout ),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hFFFE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(read_latency_shift_reg_03),
	.datab(out_valid1),
	.datac(out_data_buffer_21),
	.datad(av_readdata_pre_21),
	.cin(gnd),
	.combout(\src_payload~15_combout ),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hFFFE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(read_latency_shift_reg_03),
	.datab(out_valid1),
	.datac(out_data_buffer_20),
	.datad(av_readdata_pre_20),
	.cin(gnd),
	.combout(\src_payload~17_combout ),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hFFFE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(read_latency_shift_reg_03),
	.datab(out_valid1),
	.datac(out_data_buffer_19),
	.datad(av_readdata_pre_19),
	.cin(gnd),
	.combout(\src_payload~19_combout ),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hFFFE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~29 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_27),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\src_data[2]~29_combout ),
	.cout());
defparam \src_data[2]~29 .lut_mask = 16'hFFFE;
defparam \src_data[2]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~38 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_44),
	.datad(av_readdata_pre_45),
	.cin(gnd),
	.combout(\src_data[4]~38_combout ),
	.cout());
defparam \src_data[4]~38 .lut_mask = 16'hFFFE;
defparam \src_data[4]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~42 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_54),
	.datad(av_readdata_pre_55),
	.cin(gnd),
	.combout(\src_data[5]~42_combout ),
	.cout());
defparam \src_data[5]~42 .lut_mask = 16'hFFFE;
defparam \src_data[5]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~46 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_64),
	.datad(av_readdata_pre_65),
	.cin(gnd),
	.combout(\src_data[6]~46_combout ),
	.cout());
defparam \src_data[6]~46 .lut_mask = 16'hFFFE;
defparam \src_data[6]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~50 (
	.dataa(read_latency_shift_reg_01),
	.datab(read_latency_shift_reg_07),
	.datac(av_readdata_pre_74),
	.datad(av_readdata_pre_75),
	.cin(gnd),
	.combout(\src_data[7]~50_combout ),
	.cout());
defparam \src_data[7]~50 .lut_mask = 16'hFFFE;
defparam \src_data[7]~50 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_0_rsp_mux_001 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	read_latency_shift_reg_01,
	mem_86_01,
	mem_68_01,
	src1_valid,
	src_payload,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	src_payload1,
	WideOr1,
	out_data_buffer_3,
	src_payload2,
	out_data_buffer_16,
	src_payload3,
	out_data_buffer_20,
	src_payload4,
	out_data_buffer_21,
	src_payload5)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
input 	read_latency_shift_reg_01;
input 	mem_86_01;
input 	mem_68_01;
input 	src1_valid;
output 	src_payload;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid;
output 	src_payload1;
output 	WideOr1;
input 	out_data_buffer_3;
output 	src_payload2;
input 	out_data_buffer_16;
output 	src_payload3;
input 	out_data_buffer_20;
output 	src_payload4;
input 	out_data_buffer_21;
output 	src_payload5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_86_01),
	.datac(mem_68_01),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hFEFE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hFEFE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(src1_valid),
	.datab(src_payload),
	.datac(out_valid),
	.datad(src_payload1),
	.cin(gnd),
	.combout(WideOr1),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(out_data_buffer_3),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hAFFA;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(out_data_buffer_16),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hAFFA;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(out_data_buffer_20),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hAFFA;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(out_data_buffer_21),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hAFFA;
defparam \src_payload~5 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_mm_interconnect_1 (
	wire_pll7_clk_1,
	altera_reset_synchronizer_int_chain_out,
	out_valid,
	m0_read,
	CY7C67200_IF_0_hpi_read,
	out_payload_37,
	CY7C67200_IF_0_hpi_write,
	waitrequest_reset_override,
	av_waitrequest_generated,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	oDATA_0,
	oDATA_1,
	oDATA_2,
	oDATA_3,
	oDATA_4,
	oDATA_5,
	oDATA_6,
	oDATA_7,
	oDATA_8,
	oDATA_9,
	oDATA_10,
	oDATA_11,
	oDATA_12,
	oDATA_13,
	oDATA_14,
	oDATA_15,
	av_begintransfer)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	out_valid;
input 	m0_read;
output 	CY7C67200_IF_0_hpi_read;
input 	out_payload_37;
output 	CY7C67200_IF_0_hpi_write;
output 	waitrequest_reset_override;
output 	av_waitrequest_generated;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
input 	oDATA_0;
input 	oDATA_1;
input 	oDATA_2;
input 	oDATA_3;
input 	oDATA_4;
input 	oDATA_5;
input 	oDATA_6;
input 	oDATA_7;
input 	oDATA_8;
input 	oDATA_9;
input 	oDATA_10;
input 	oDATA_11;
input 	oDATA_12;
input 	oDATA_13;
input 	oDATA_14;
input 	oDATA_15;
output 	av_begintransfer;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



usb_system_altera_merlin_slave_translator_10 cy7c67200_if_0_hpi_translator(
	.clk(wire_pll7_clk_1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid),
	.m0_read(m0_read),
	.av_read(CY7C67200_IF_0_hpi_read),
	.out_payload_37(out_payload_37),
	.av_write(CY7C67200_IF_0_hpi_write),
	.waitrequest_reset_override1(waitrequest_reset_override),
	.av_waitrequest_generated(av_waitrequest_generated),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,oDATA_15,oDATA_14,oDATA_13,oDATA_12,oDATA_11,oDATA_10,oDATA_9,oDATA_8,oDATA_7,oDATA_6,oDATA_5,oDATA_4,oDATA_3,oDATA_2,oDATA_1,oDATA_0}),
	.av_begintransfer(av_begintransfer));

endmodule

module usb_system_altera_merlin_slave_translator_10 (
	clk,
	reset,
	out_valid,
	m0_read,
	av_read,
	out_payload_37,
	av_write,
	waitrequest_reset_override1,
	av_waitrequest_generated,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata,
	av_begintransfer)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	out_valid;
input 	m0_read;
output 	av_read;
input 	out_payload_37;
output 	av_write;
output 	waitrequest_reset_override1;
output 	av_waitrequest_generated;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
input 	[31:0] av_readdata;
output 	av_begintransfer;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_waitrequest_generated~0_combout ;
wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter[1]~q ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter[2]~q ;
wire \read_latency_shift_reg~0_combout ;


cycloneive_lcell_comb \av_read~0 (
	.dataa(m0_read),
	.datab(\wait_latency_counter[2]~q ),
	.datac(\wait_latency_counter[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_read),
	.cout());
defparam \av_read~0 .lut_mask = 16'hFEFE;
defparam \av_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_write~0 (
	.dataa(\av_waitrequest_generated~0_combout ),
	.datab(\wait_latency_counter[1]~q ),
	.datac(\wait_latency_counter[0]~q ),
	.datad(\wait_latency_counter[2]~q ),
	.cin(gnd),
	.combout(av_write),
	.cout());
defparam \av_write~0 .lut_mask = 16'hBFEF;
defparam \av_write~0 .sum_lutc_input = "datac";

dffeas waitrequest_reset_override(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_reset_override1),
	.prn(vcc));
defparam waitrequest_reset_override.is_wysiwyg = "true";
defparam waitrequest_reset_override.power_up = "low";

cycloneive_lcell_comb \av_waitrequest_generated~1 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(\wait_latency_counter[1]~q ),
	.datac(\av_waitrequest_generated~0_combout ),
	.datad(\wait_latency_counter[2]~q ),
	.cin(gnd),
	.combout(av_waitrequest_generated),
	.cout());
defparam \av_waitrequest_generated~1 .lut_mask = 16'hBEFF;
defparam \av_waitrequest_generated~1 .sum_lutc_input = "datac";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

cycloneive_lcell_comb \av_begintransfer~2 (
	.dataa(out_valid),
	.datab(out_payload_37),
	.datac(m0_read),
	.datad(gnd),
	.cin(gnd),
	.combout(av_begintransfer),
	.cout());
defparam \av_begintransfer~2 .lut_mask = 16'hFEFE;
defparam \av_begintransfer~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest_generated~0 (
	.dataa(out_valid),
	.datab(out_payload_37),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest_generated~0_combout ),
	.cout());
defparam \av_waitrequest_generated~0 .lut_mask = 16'hEEEE;
defparam \av_waitrequest_generated~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~0 (
	.dataa(waitrequest_reset_override1),
	.datab(av_waitrequest_generated),
	.datac(m0_read),
	.datad(\av_waitrequest_generated~0_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.cout());
defparam \wait_latency_counter~0 .lut_mask = 16'hFFFE;
defparam \wait_latency_counter~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(av_begintransfer),
	.datac(waitrequest_reset_override1),
	.datad(av_waitrequest_generated),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFFFD;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter~0_combout ),
	.datab(gnd),
	.datac(\wait_latency_counter[1]~q ),
	.datad(\wait_latency_counter[0]~q ),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[1]~q ),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter~1 (
	.dataa(\wait_latency_counter~0_combout ),
	.datab(\wait_latency_counter[2]~q ),
	.datac(\wait_latency_counter[1]~q ),
	.datad(\wait_latency_counter[0]~q ),
	.cin(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.cout());
defparam \wait_latency_counter~1 .lut_mask = 16'hEBBE;
defparam \wait_latency_counter~1 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[2] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[2]~q ),
	.prn(vcc));
defparam \wait_latency_counter[2] .is_wysiwyg = "true";
defparam \wait_latency_counter[2] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(av_waitrequest_generated),
	.datab(gnd),
	.datac(m0_read),
	.datad(waitrequest_reset_override1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFF5;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_red_leds (
	W_alu_result_7,
	W_alu_result_4,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	writedata,
	Equal3,
	always0,
	reset_n,
	mem_used_1,
	always01,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_4;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_16;
output 	data_out_17;
input 	[31:0] writedata;
input 	Equal3;
input 	always0;
input 	reset_n;
input 	mem_used_1;
output 	always01;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~2_combout ;
wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(writedata[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(writedata[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

cycloneive_lcell_comb \always0~1 (
	.dataa(W_alu_result_5),
	.datab(mem_used_1),
	.datac(Equal3),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(always01),
	.cout());
defparam \always0~1 .lut_mask = 16'hFFF7;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAFFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAFFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAFFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAFFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAFFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAFFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAFFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAFFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[8] (
	.dataa(data_out_8),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_8),
	.cout());
defparam \readdata[8] .lut_mask = 16'hAFFF;
defparam \readdata[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[9] (
	.dataa(data_out_9),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_9),
	.cout());
defparam \readdata[9] .lut_mask = 16'hAFFF;
defparam \readdata[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[10] (
	.dataa(data_out_10),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_10),
	.cout());
defparam \readdata[10] .lut_mask = 16'hAFFF;
defparam \readdata[10] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[11] (
	.dataa(data_out_11),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_11),
	.cout());
defparam \readdata[11] .lut_mask = 16'hAFFF;
defparam \readdata[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[12] (
	.dataa(data_out_12),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_12),
	.cout());
defparam \readdata[12] .lut_mask = 16'hAFFF;
defparam \readdata[12] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[13] (
	.dataa(data_out_13),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_13),
	.cout());
defparam \readdata[13] .lut_mask = 16'hAFFF;
defparam \readdata[13] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[14] (
	.dataa(data_out_14),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_14),
	.cout());
defparam \readdata[14] .lut_mask = 16'hAFFF;
defparam \readdata[14] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[15] (
	.dataa(data_out_15),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_15),
	.cout());
defparam \readdata[15] .lut_mask = 16'hAFFF;
defparam \readdata[15] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[16] (
	.dataa(data_out_16),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_16),
	.cout());
defparam \readdata[16] .lut_mask = 16'hAFFF;
defparam \readdata[16] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[17] (
	.dataa(data_out_17),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_17),
	.cout());
defparam \readdata[17] .lut_mask = 16'hAFFF;
defparam \readdata[17] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~2 (
	.dataa(always0),
	.datab(always01),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hEFFF;
defparam \always0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hBBBB;
defparam \always0~0 .sum_lutc_input = "datac";

endmodule

module usb_system_usb_system_sdram (
	wire_pll7_clk_0,
	m_addr_0,
	m_addr_1,
	m_addr_2,
	m_addr_3,
	m_addr_4,
	m_addr_5,
	m_addr_6,
	m_addr_7,
	m_addr_8,
	m_addr_9,
	oe1,
	m_addr_10,
	m_addr_11,
	m_addr_12,
	m_bank_0,
	m_bank_1,
	m_cmd_1,
	m_cmd_3,
	m_dqm_0,
	m_dqm_1,
	m_dqm_2,
	m_dqm_3,
	m_cmd_2,
	m_cmd_0,
	entries_1,
	entries_0,
	altera_reset_synchronizer_int_chain_out,
	last_cycle,
	saved_grant_1,
	WideOr1,
	src_payload,
	src_data_68,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	src_data_61,
	src_data_60,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	out_data_buffer_32,
	out_data_buffer_321,
	out_data_buffer_33,
	out_data_buffer_331,
	out_data_buffer_34,
	out_data_buffer_341,
	out_data_buffer_35,
	out_data_buffer_351,
	m_data_0,
	m_data_1,
	m_data_2,
	m_data_3,
	m_data_4,
	m_data_5,
	m_data_6,
	m_data_7,
	m_data_8,
	m_data_9,
	m_data_10,
	m_data_11,
	m_data_12,
	m_data_13,
	m_data_14,
	m_data_15,
	m_data_16,
	m_data_17,
	m_data_18,
	m_data_19,
	m_data_20,
	m_data_21,
	m_data_22,
	m_data_23,
	m_data_24,
	m_data_25,
	m_data_26,
	m_data_27,
	m_data_28,
	m_data_29,
	m_data_30,
	m_data_31,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	za_valid1,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_22,
	za_data_23,
	za_data_24,
	za_data_25,
	za_data_26,
	za_data_11,
	za_data_13,
	za_data_16,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_10,
	za_data_9,
	za_data_8,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_18,
	za_data_19,
	za_data_17,
	za_data_21,
	za_data_27,
	za_data_28,
	za_data_31,
	za_data_30,
	za_data_29,
	m0_write,
	sdram_wire_dq_0,
	sdram_wire_dq_1,
	sdram_wire_dq_2,
	sdram_wire_dq_3,
	sdram_wire_dq_4,
	sdram_wire_dq_5,
	sdram_wire_dq_6,
	sdram_wire_dq_7,
	sdram_wire_dq_8,
	sdram_wire_dq_9,
	sdram_wire_dq_10,
	sdram_wire_dq_11,
	sdram_wire_dq_12,
	sdram_wire_dq_13,
	sdram_wire_dq_14,
	sdram_wire_dq_15,
	sdram_wire_dq_16,
	sdram_wire_dq_17,
	sdram_wire_dq_18,
	sdram_wire_dq_19,
	sdram_wire_dq_20,
	sdram_wire_dq_21,
	sdram_wire_dq_22,
	sdram_wire_dq_23,
	sdram_wire_dq_24,
	sdram_wire_dq_25,
	sdram_wire_dq_26,
	sdram_wire_dq_27,
	sdram_wire_dq_28,
	sdram_wire_dq_29,
	sdram_wire_dq_30,
	sdram_wire_dq_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	m_addr_0;
output 	m_addr_1;
output 	m_addr_2;
output 	m_addr_3;
output 	m_addr_4;
output 	m_addr_5;
output 	m_addr_6;
output 	m_addr_7;
output 	m_addr_8;
output 	m_addr_9;
output 	oe1;
output 	m_addr_10;
output 	m_addr_11;
output 	m_addr_12;
output 	m_bank_0;
output 	m_bank_1;
output 	m_cmd_1;
output 	m_cmd_3;
output 	m_dqm_0;
output 	m_dqm_1;
output 	m_dqm_2;
output 	m_dqm_3;
output 	m_cmd_2;
output 	m_cmd_0;
output 	entries_1;
output 	entries_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	last_cycle;
input 	saved_grant_1;
input 	WideOr1;
input 	src_payload;
input 	src_data_68;
input 	src_data_48;
input 	src_data_62;
input 	src_data_49;
input 	src_data_51;
input 	src_data_50;
input 	src_data_53;
input 	src_data_52;
input 	src_data_55;
input 	src_data_54;
input 	src_data_57;
input 	src_data_56;
input 	src_data_59;
input 	src_data_58;
input 	src_data_61;
input 	src_data_60;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	out_data_buffer_32;
input 	out_data_buffer_321;
input 	out_data_buffer_33;
input 	out_data_buffer_331;
input 	out_data_buffer_34;
input 	out_data_buffer_341;
input 	out_data_buffer_35;
input 	out_data_buffer_351;
output 	m_data_0;
output 	m_data_1;
output 	m_data_2;
output 	m_data_3;
output 	m_data_4;
output 	m_data_5;
output 	m_data_6;
output 	m_data_7;
output 	m_data_8;
output 	m_data_9;
output 	m_data_10;
output 	m_data_11;
output 	m_data_12;
output 	m_data_13;
output 	m_data_14;
output 	m_data_15;
output 	m_data_16;
output 	m_data_17;
output 	m_data_18;
output 	m_data_19;
output 	m_data_20;
output 	m_data_21;
output 	m_data_22;
output 	m_data_23;
output 	m_data_24;
output 	m_data_25;
output 	m_data_26;
output 	m_data_27;
output 	m_data_28;
output 	m_data_29;
output 	m_data_30;
output 	m_data_31;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
output 	za_valid1;
output 	za_data_0;
output 	za_data_1;
output 	za_data_2;
output 	za_data_3;
output 	za_data_4;
output 	za_data_22;
output 	za_data_23;
output 	za_data_24;
output 	za_data_25;
output 	za_data_26;
output 	za_data_11;
output 	za_data_13;
output 	za_data_16;
output 	za_data_12;
output 	za_data_5;
output 	za_data_14;
output 	za_data_15;
output 	za_data_10;
output 	za_data_9;
output 	za_data_8;
output 	za_data_7;
output 	za_data_6;
output 	za_data_20;
output 	za_data_18;
output 	za_data_19;
output 	za_data_17;
output 	za_data_21;
output 	za_data_27;
output 	za_data_28;
output 	za_data_31;
output 	za_data_30;
output 	za_data_29;
input 	m0_write;
input 	sdram_wire_dq_0;
input 	sdram_wire_dq_1;
input 	sdram_wire_dq_2;
input 	sdram_wire_dq_3;
input 	sdram_wire_dq_4;
input 	sdram_wire_dq_5;
input 	sdram_wire_dq_6;
input 	sdram_wire_dq_7;
input 	sdram_wire_dq_8;
input 	sdram_wire_dq_9;
input 	sdram_wire_dq_10;
input 	sdram_wire_dq_11;
input 	sdram_wire_dq_12;
input 	sdram_wire_dq_13;
input 	sdram_wire_dq_14;
input 	sdram_wire_dq_15;
input 	sdram_wire_dq_16;
input 	sdram_wire_dq_17;
input 	sdram_wire_dq_18;
input 	sdram_wire_dq_19;
input 	sdram_wire_dq_20;
input 	sdram_wire_dq_21;
input 	sdram_wire_dq_22;
input 	sdram_wire_dq_23;
input 	sdram_wire_dq_24;
input 	sdram_wire_dq_25;
input 	sdram_wire_dq_26;
input 	sdram_wire_dq_27;
input 	sdram_wire_dq_28;
input 	sdram_wire_dq_29;
input 	sdram_wire_dq_30;
input 	sdram_wire_dq_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_usb_system_sdram_input_efifo_module|Equal1~0_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[46]~0_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[61]~1_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[60]~2_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[47]~3_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[49]~4_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[48]~5_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[51]~6_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[50]~7_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[53]~8_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[52]~9_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[55]~10_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[54]~11_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[57]~12_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[56]~13_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[59]~14_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[58]~15_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[36]~16_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[37]~17_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[38]~18_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[39]~19_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[40]~20_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[41]~21_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[42]~22_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[43]~23_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[44]~24_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[45]~25_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[32]~26_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[33]~27_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[34]~28_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[35]~29_combout ;
wire \comb~0_combout ;
wire \comb~1_combout ;
wire \comb~2_combout ;
wire \comb~3_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[0]~30_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[1]~31_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[2]~32_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[3]~33_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[4]~34_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[5]~35_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[6]~36_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[7]~37_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[8]~38_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[9]~39_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[10]~40_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[11]~41_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[12]~42_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[13]~43_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[14]~44_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[15]~45_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[16]~46_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[17]~47_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[18]~48_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[19]~49_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[20]~50_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[21]~51_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[22]~52_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[23]~53_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[24]~54_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[25]~55_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[26]~56_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[27]~57_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[28]~58_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[29]~59_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[30]~60_combout ;
wire \the_usb_system_sdram_input_efifo_module|rd_data[31]~61_combout ;
wire \Add0~0_combout ;
wire \refresh_counter~9_combout ;
wire \refresh_counter[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \refresh_counter[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \refresh_counter[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \refresh_counter~8_combout ;
wire \refresh_counter[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \refresh_counter~6_combout ;
wire \refresh_counter[4]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \refresh_counter~7_combout ;
wire \refresh_counter[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \refresh_counter~5_combout ;
wire \refresh_counter[6]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \refresh_counter[7]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \refresh_counter[8]~13_combout ;
wire \refresh_counter[8]~q ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \refresh_counter~4_combout ;
wire \refresh_counter[9]~q ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \refresh_counter~1_combout ;
wire \refresh_counter[10]~q ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \refresh_counter~3_combout ;
wire \refresh_counter[11]~q ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \refresh_counter~2_combout ;
wire \refresh_counter[12]~q ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \refresh_counter~0_combout ;
wire \refresh_counter[13]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \i_next.000~0_combout ;
wire \i_next.000~q ;
wire \Selector7~0_combout ;
wire \i_state.000~q ;
wire \Selector18~0_combout ;
wire \Selector8~0_combout ;
wire \i_state.001~q ;
wire \Selector16~0_combout ;
wire \Selector6~0_combout ;
wire \i_refs[0]~q ;
wire \Selector5~0_combout ;
wire \i_refs[1]~q ;
wire \Selector4~0_combout ;
wire \Selector4~1_combout ;
wire \i_refs[2]~q ;
wire \Selector18~1_combout ;
wire \Selector16~1_combout ;
wire \i_next.010~q ;
wire \i_count[0]~4_combout ;
wire \i_count[0]~1_combout ;
wire \i_count[0]~5_combout ;
wire \i_count[0]~q ;
wire \i_count[1]~2_combout ;
wire \i_count[1]~3_combout ;
wire \i_count[1]~q ;
wire \Selector13~0_combout ;
wire \Selector13~1_combout ;
wire \i_count[2]~q ;
wire \Selector9~0_combout ;
wire \i_state.010~q ;
wire \Selector18~2_combout ;
wire \i_next.111~q ;
wire \Selector12~0_combout ;
wire \i_state.111~q ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \i_state.011~q ;
wire \i_count[0]~0_combout ;
wire \WideOr6~0_combout ;
wire \Selector17~0_combout ;
wire \i_next.101~q ;
wire \i_state.101~0_combout ;
wire \i_state.101~q ;
wire \init_done~0_combout ;
wire \init_done~q ;
wire \Selector24~1_combout ;
wire \Selector32~0_combout ;
wire \active_rnw~q ;
wire \Selector25~5_combout ;
wire \Selector25~6_combout ;
wire \m_state.000000010~q ;
wire \active_addr[10]~q ;
wire \pending~0_combout ;
wire \active_addr[24]~q ;
wire \pending~1_combout ;
wire \active_addr[12]~q ;
wire \active_addr[13]~q ;
wire \pending~2_combout ;
wire \active_addr[14]~q ;
wire \active_addr[15]~q ;
wire \pending~3_combout ;
wire \pending~4_combout ;
wire \active_addr[16]~q ;
wire \active_addr[17]~q ;
wire \pending~5_combout ;
wire \active_addr[18]~q ;
wire \active_addr[19]~q ;
wire \pending~6_combout ;
wire \active_addr[20]~q ;
wire \active_addr[21]~q ;
wire \pending~7_combout ;
wire \active_addr[22]~q ;
wire \active_addr[23]~q ;
wire \pending~8_combout ;
wire \pending~9_combout ;
wire \pending~10_combout ;
wire \m_next~22_combout ;
wire \Selector25~4_combout ;
wire \Selector38~0_combout ;
wire \m_next~21_combout ;
wire \Selector29~0_combout ;
wire \Selector39~1_combout ;
wire \Selector39~2_combout ;
wire \Selector39~3_combout ;
wire \WideOr10~0_combout ;
wire \Selector27~0_combout ;
wire \Selector35~5_combout ;
wire \Selector34~1_combout ;
wire \Selector35~3_combout ;
wire \Selector35~4_combout ;
wire \Selector34~2_combout ;
wire \m_next.000010000~q ;
wire \Selector27~1_combout ;
wire \Selector28~0_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \WideOr8~0_combout ;
wire \Selector27~5_combout ;
wire \Selector27~6_combout ;
wire \m_state.000010000~q ;
wire \Selector39~0_combout ;
wire \Selector39~4_combout ;
wire \Selector39~5_combout ;
wire \m_count[0]~q ;
wire \Selector38~1_combout ;
wire \Selector38~2_combout ;
wire \Selector38~3_combout ;
wire \Selector38~4_combout ;
wire \m_count[1]~q ;
wire \Selector29~1_combout ;
wire \m_state.000100000~q ;
wire \Selector30~0_combout ;
wire \Selector30~1_combout ;
wire \m_state.001000000~q ;
wire \Selector33~0_combout ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \m_next.010000000~q ;
wire \Selector31~0_combout ;
wire \m_state.010000000~q ;
wire \Selector35~2_combout ;
wire \Selector34~0_combout ;
wire \m_next.000001000~q ;
wire \Selector27~2_combout ;
wire \m_state.000001000~q ;
wire \WideOr9~0_combout ;
wire \Selector32~1_combout ;
wire \m_state.100000000~q ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector26~2_combout ;
wire \m_state.000000100~q ;
wire \Selector24~0_combout ;
wire \Selector35~6_combout ;
wire \Selector33~1_combout ;
wire \Selector33~2_combout ;
wire \Selector33~3_combout ;
wire \Selector33~4_combout ;
wire \m_next.000000001~q ;
wire \Selector24~2_combout ;
wire \m_state.000000001~q ;
wire \Selector23~0_combout ;
wire \ack_refresh_request~q ;
wire \refresh_request~0_combout ;
wire \refresh_request~q ;
wire \active_cs_n~0_combout ;
wire \active_cs_n~1_combout ;
wire \active_cs_n~q ;
wire \pending~combout ;
wire \active_rnw~2_combout ;
wire \active_rnw~4_combout ;
wire \active_rnw~3_combout ;
wire \active_addr[11]~q ;
wire \Selector41~0_combout ;
wire \Selector41~1_combout ;
wire \f_pop~q ;
wire \m_addr[3]~0_combout ;
wire \active_addr[0]~q ;
wire \i_addr[12]~q ;
wire \Selector116~0_combout ;
wire \Selector116~1_combout ;
wire \m_addr[3]~1_combout ;
wire \m_addr[3]~2_combout ;
wire \active_addr[1]~q ;
wire \Selector115~0_combout ;
wire \Selector115~1_combout ;
wire \active_addr[2]~q ;
wire \Selector114~0_combout ;
wire \Selector114~1_combout ;
wire \active_addr[3]~q ;
wire \Selector113~0_combout ;
wire \Selector113~1_combout ;
wire \active_addr[4]~q ;
wire \f_select~combout ;
wire \Selector112~0_combout ;
wire \Selector112~1_combout ;
wire \active_addr[5]~q ;
wire \Selector111~0_combout ;
wire \Selector111~1_combout ;
wire \active_addr[6]~q ;
wire \Selector110~0_combout ;
wire \Selector110~1_combout ;
wire \active_addr[7]~q ;
wire \Selector109~0_combout ;
wire \Selector109~1_combout ;
wire \active_addr[8]~q ;
wire \Selector108~0_combout ;
wire \Selector108~1_combout ;
wire \active_addr[9]~q ;
wire \Selector107~0_combout ;
wire \Selector107~1_combout ;
wire \always5~0_combout ;
wire \Selector106~2_combout ;
wire \Selector106~3_combout ;
wire \Selector105~2_combout ;
wire \Selector105~3_combout ;
wire \Selector104~2_combout ;
wire \Selector104~3_combout ;
wire \Selector118~0_combout ;
wire \WideOr16~0_combout ;
wire \Selector117~0_combout ;
wire \Selector2~0_combout ;
wire \i_cmd[1]~q ;
wire \Selector21~0_combout ;
wire \Selector21~1_combout ;
wire \Selector0~0_combout ;
wire \i_cmd[3]~q ;
wire \Selector19~0_combout ;
wire \Selector19~1_combout ;
wire \Selector19~2_combout ;
wire \Selector19~3_combout ;
wire \active_dqm[0]~q ;
wire \Selector154~0_combout ;
wire \active_dqm[1]~q ;
wire \Selector153~0_combout ;
wire \active_dqm[2]~q ;
wire \Selector152~0_combout ;
wire \active_dqm[3]~q ;
wire \Selector151~0_combout ;
wire \Selector1~0_combout ;
wire \i_cmd[2]~q ;
wire \Selector20~0_combout ;
wire \Selector3~0_combout ;
wire \i_cmd[0]~q ;
wire \Selector22~0_combout ;
wire \Selector22~1_combout ;
wire \active_data[0]~q ;
wire \Selector150~0_combout ;
wire \m_data[30]~0_combout ;
wire \Selector150~1_combout ;
wire \active_data[1]~q ;
wire \Selector149~0_combout ;
wire \Selector149~1_combout ;
wire \active_data[2]~q ;
wire \Selector148~0_combout ;
wire \Selector148~1_combout ;
wire \active_data[3]~q ;
wire \Selector147~0_combout ;
wire \Selector147~1_combout ;
wire \active_data[4]~q ;
wire \Selector146~0_combout ;
wire \Selector146~1_combout ;
wire \active_data[5]~q ;
wire \Selector145~0_combout ;
wire \Selector145~1_combout ;
wire \active_data[6]~q ;
wire \Selector144~0_combout ;
wire \Selector144~1_combout ;
wire \active_data[7]~q ;
wire \Selector143~0_combout ;
wire \Selector143~1_combout ;
wire \active_data[8]~q ;
wire \Selector142~0_combout ;
wire \Selector142~1_combout ;
wire \active_data[9]~q ;
wire \Selector141~0_combout ;
wire \Selector141~1_combout ;
wire \active_data[10]~q ;
wire \Selector140~0_combout ;
wire \Selector140~1_combout ;
wire \active_data[11]~q ;
wire \Selector139~0_combout ;
wire \Selector139~1_combout ;
wire \active_data[12]~q ;
wire \Selector138~0_combout ;
wire \Selector138~1_combout ;
wire \active_data[13]~q ;
wire \Selector137~0_combout ;
wire \Selector137~1_combout ;
wire \active_data[14]~q ;
wire \Selector136~0_combout ;
wire \Selector136~1_combout ;
wire \active_data[15]~q ;
wire \Selector135~0_combout ;
wire \Selector135~1_combout ;
wire \active_data[16]~q ;
wire \Selector134~0_combout ;
wire \Selector134~1_combout ;
wire \active_data[17]~q ;
wire \Selector133~0_combout ;
wire \Selector133~1_combout ;
wire \active_data[18]~q ;
wire \Selector132~0_combout ;
wire \Selector132~1_combout ;
wire \active_data[19]~q ;
wire \Selector131~0_combout ;
wire \Selector131~1_combout ;
wire \active_data[20]~q ;
wire \Selector130~0_combout ;
wire \Selector130~1_combout ;
wire \active_data[21]~q ;
wire \Selector129~0_combout ;
wire \Selector129~1_combout ;
wire \active_data[22]~q ;
wire \Selector128~0_combout ;
wire \Selector128~1_combout ;
wire \active_data[23]~q ;
wire \Selector127~0_combout ;
wire \Selector127~1_combout ;
wire \active_data[24]~q ;
wire \Selector126~0_combout ;
wire \Selector126~1_combout ;
wire \active_data[25]~q ;
wire \Selector125~0_combout ;
wire \Selector125~1_combout ;
wire \active_data[26]~q ;
wire \Selector124~0_combout ;
wire \Selector124~1_combout ;
wire \active_data[27]~q ;
wire \Selector123~0_combout ;
wire \Selector123~1_combout ;
wire \active_data[28]~q ;
wire \Selector122~0_combout ;
wire \Selector122~1_combout ;
wire \active_data[29]~q ;
wire \Selector121~0_combout ;
wire \Selector121~1_combout ;
wire \active_data[30]~q ;
wire \Selector120~0_combout ;
wire \Selector120~1_combout ;
wire \active_data[31]~q ;
wire \Selector119~0_combout ;
wire \Selector119~1_combout ;
wire \Equal4~0_combout ;
wire \rd_valid[0]~q ;
wire \rd_valid[1]~q ;
wire \rd_valid[2]~q ;


usb_system_usb_system_sdram_input_efifo_module the_usb_system_sdram_input_efifo_module(
	.clk(wire_pll7_clk_0),
	.f_pop(\f_pop~q ),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.Equal1(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.rd_data_46(\the_usb_system_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.rd_data_61(\the_usb_system_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.rd_data_60(\the_usb_system_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.rd_data_47(\the_usb_system_sdram_input_efifo_module|rd_data[47]~3_combout ),
	.rd_data_49(\the_usb_system_sdram_input_efifo_module|rd_data[49]~4_combout ),
	.rd_data_48(\the_usb_system_sdram_input_efifo_module|rd_data[48]~5_combout ),
	.rd_data_51(\the_usb_system_sdram_input_efifo_module|rd_data[51]~6_combout ),
	.rd_data_50(\the_usb_system_sdram_input_efifo_module|rd_data[50]~7_combout ),
	.rd_data_53(\the_usb_system_sdram_input_efifo_module|rd_data[53]~8_combout ),
	.rd_data_52(\the_usb_system_sdram_input_efifo_module|rd_data[52]~9_combout ),
	.rd_data_55(\the_usb_system_sdram_input_efifo_module|rd_data[55]~10_combout ),
	.rd_data_54(\the_usb_system_sdram_input_efifo_module|rd_data[54]~11_combout ),
	.rd_data_57(\the_usb_system_sdram_input_efifo_module|rd_data[57]~12_combout ),
	.rd_data_56(\the_usb_system_sdram_input_efifo_module|rd_data[56]~13_combout ),
	.rd_data_59(\the_usb_system_sdram_input_efifo_module|rd_data[59]~14_combout ),
	.rd_data_58(\the_usb_system_sdram_input_efifo_module|rd_data[58]~15_combout ),
	.pending(\pending~combout ),
	.rd_data_36(\the_usb_system_sdram_input_efifo_module|rd_data[36]~16_combout ),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.rd_data_37(\the_usb_system_sdram_input_efifo_module|rd_data[37]~17_combout ),
	.rd_data_38(\the_usb_system_sdram_input_efifo_module|rd_data[38]~18_combout ),
	.rd_data_39(\the_usb_system_sdram_input_efifo_module|rd_data[39]~19_combout ),
	.rd_data_40(\the_usb_system_sdram_input_efifo_module|rd_data[40]~20_combout ),
	.f_select(\f_select~combout ),
	.rd_data_41(\the_usb_system_sdram_input_efifo_module|rd_data[41]~21_combout ),
	.rd_data_42(\the_usb_system_sdram_input_efifo_module|rd_data[42]~22_combout ),
	.rd_data_43(\the_usb_system_sdram_input_efifo_module|rd_data[43]~23_combout ),
	.rd_data_44(\the_usb_system_sdram_input_efifo_module|rd_data[44]~24_combout ),
	.rd_data_45(\the_usb_system_sdram_input_efifo_module|rd_data[45]~25_combout ),
	.rd_data_32(\the_usb_system_sdram_input_efifo_module|rd_data[32]~26_combout ),
	.rd_data_33(\the_usb_system_sdram_input_efifo_module|rd_data[33]~27_combout ),
	.rd_data_34(\the_usb_system_sdram_input_efifo_module|rd_data[34]~28_combout ),
	.rd_data_35(\the_usb_system_sdram_input_efifo_module|rd_data[35]~29_combout ),
	.last_cycle(last_cycle),
	.WideOr1(WideOr1),
	.src_payload(src_payload),
	.src_data_68(src_data_68),
	.src_data_48(src_data_48),
	.src_data_62(src_data_62),
	.src_data_49(src_data_49),
	.src_data_51(src_data_51),
	.src_data_50(src_data_50),
	.src_data_53(src_data_53),
	.src_data_52(src_data_52),
	.src_data_55(src_data_55),
	.src_data_54(src_data_54),
	.src_data_57(src_data_57),
	.src_data_56(src_data_56),
	.src_data_59(src_data_59),
	.src_data_58(src_data_58),
	.src_data_61(src_data_61),
	.src_data_60(src_data_60),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_46),
	.src_data_47(src_data_47),
	.comb(\comb~0_combout ),
	.comb1(\comb~1_combout ),
	.comb2(\comb~2_combout ),
	.comb3(\comb~3_combout ),
	.rd_data_0(\the_usb_system_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.rd_data_1(\the_usb_system_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.rd_data_2(\the_usb_system_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.rd_data_3(\the_usb_system_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.rd_data_4(\the_usb_system_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.rd_data_5(\the_usb_system_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.rd_data_6(\the_usb_system_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.rd_data_7(\the_usb_system_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.rd_data_8(\the_usb_system_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.rd_data_9(\the_usb_system_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.rd_data_10(\the_usb_system_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.rd_data_11(\the_usb_system_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.rd_data_12(\the_usb_system_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.rd_data_13(\the_usb_system_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.rd_data_14(\the_usb_system_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.rd_data_15(\the_usb_system_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.rd_data_16(\the_usb_system_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.rd_data_17(\the_usb_system_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.rd_data_18(\the_usb_system_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.rd_data_19(\the_usb_system_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.rd_data_20(\the_usb_system_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.rd_data_21(\the_usb_system_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.rd_data_22(\the_usb_system_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.rd_data_23(\the_usb_system_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.rd_data_24(\the_usb_system_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.rd_data_25(\the_usb_system_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.rd_data_26(\the_usb_system_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.rd_data_27(\the_usb_system_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.rd_data_28(\the_usb_system_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.rd_data_29(\the_usb_system_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.rd_data_30(\the_usb_system_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.rd_data_31(\the_usb_system_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.m0_write(m0_write));

cycloneive_lcell_comb \comb~0 (
	.dataa(out_data_buffer_32),
	.datab(saved_grant_1),
	.datac(out_data_buffer_321),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'h7FFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~1 (
	.dataa(out_data_buffer_33),
	.datab(saved_grant_1),
	.datac(out_data_buffer_331),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'h7FFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~2 (
	.dataa(out_data_buffer_34),
	.datab(saved_grant_1),
	.datac(out_data_buffer_341),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
defparam \comb~2 .lut_mask = 16'h7FFF;
defparam \comb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~3 (
	.dataa(out_data_buffer_35),
	.datab(saved_grant_1),
	.datac(out_data_buffer_351),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~3_combout ),
	.cout());
defparam \comb~3 .lut_mask = 16'h7FFF;
defparam \comb~3 .sum_lutc_input = "datac";

dffeas \m_addr[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector116~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_0),
	.prn(vcc));
defparam \m_addr[0] .is_wysiwyg = "true";
defparam \m_addr[0] .power_up = "low";

dffeas \m_addr[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector115~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_1),
	.prn(vcc));
defparam \m_addr[1] .is_wysiwyg = "true";
defparam \m_addr[1] .power_up = "low";

dffeas \m_addr[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector114~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_2),
	.prn(vcc));
defparam \m_addr[2] .is_wysiwyg = "true";
defparam \m_addr[2] .power_up = "low";

dffeas \m_addr[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector113~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_3),
	.prn(vcc));
defparam \m_addr[3] .is_wysiwyg = "true";
defparam \m_addr[3] .power_up = "low";

dffeas \m_addr[4] (
	.clk(wire_pll7_clk_0),
	.d(\Selector112~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_4),
	.prn(vcc));
defparam \m_addr[4] .is_wysiwyg = "true";
defparam \m_addr[4] .power_up = "low";

dffeas \m_addr[5] (
	.clk(wire_pll7_clk_0),
	.d(\Selector111~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_5),
	.prn(vcc));
defparam \m_addr[5] .is_wysiwyg = "true";
defparam \m_addr[5] .power_up = "low";

dffeas \m_addr[6] (
	.clk(wire_pll7_clk_0),
	.d(\Selector110~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_6),
	.prn(vcc));
defparam \m_addr[6] .is_wysiwyg = "true";
defparam \m_addr[6] .power_up = "low";

dffeas \m_addr[7] (
	.clk(wire_pll7_clk_0),
	.d(\Selector109~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_7),
	.prn(vcc));
defparam \m_addr[7] .is_wysiwyg = "true";
defparam \m_addr[7] .power_up = "low";

dffeas \m_addr[8] (
	.clk(wire_pll7_clk_0),
	.d(\Selector108~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_8),
	.prn(vcc));
defparam \m_addr[8] .is_wysiwyg = "true";
defparam \m_addr[8] .power_up = "low";

dffeas \m_addr[9] (
	.clk(wire_pll7_clk_0),
	.d(\Selector107~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_9),
	.prn(vcc));
defparam \m_addr[9] .is_wysiwyg = "true";
defparam \m_addr[9] .power_up = "low";

dffeas oe(
	.clk(wire_pll7_clk_0),
	.d(\always5~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(!\m_state.000010000~q ),
	.sload(gnd),
	.ena(vcc),
	.q(oe1),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

dffeas \m_addr[10] (
	.clk(wire_pll7_clk_0),
	.d(\Selector106~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_10),
	.prn(vcc));
defparam \m_addr[10] .is_wysiwyg = "true";
defparam \m_addr[10] .power_up = "low";

dffeas \m_addr[11] (
	.clk(wire_pll7_clk_0),
	.d(\Selector105~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_11),
	.prn(vcc));
defparam \m_addr[11] .is_wysiwyg = "true";
defparam \m_addr[11] .power_up = "low";

dffeas \m_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\Selector104~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_12),
	.prn(vcc));
defparam \m_addr[12] .is_wysiwyg = "true";
defparam \m_addr[12] .power_up = "low";

dffeas \m_bank[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector118~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_0),
	.prn(vcc));
defparam \m_bank[0] .is_wysiwyg = "true";
defparam \m_bank[0] .power_up = "low";

dffeas \m_bank[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector117~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_1),
	.prn(vcc));
defparam \m_bank[1] .is_wysiwyg = "true";
defparam \m_bank[1] .power_up = "low";

dffeas \m_cmd[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector21~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_1),
	.prn(vcc));
defparam \m_cmd[1] .is_wysiwyg = "true";
defparam \m_cmd[1] .power_up = "low";

dffeas \m_cmd[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector19~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_3),
	.prn(vcc));
defparam \m_cmd[3] .is_wysiwyg = "true";
defparam \m_cmd[3] .power_up = "low";

dffeas \m_dqm[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector154~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_0),
	.prn(vcc));
defparam \m_dqm[0] .is_wysiwyg = "true";
defparam \m_dqm[0] .power_up = "low";

dffeas \m_dqm[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector153~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_1),
	.prn(vcc));
defparam \m_dqm[1] .is_wysiwyg = "true";
defparam \m_dqm[1] .power_up = "low";

dffeas \m_dqm[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector152~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_2),
	.prn(vcc));
defparam \m_dqm[2] .is_wysiwyg = "true";
defparam \m_dqm[2] .power_up = "low";

dffeas \m_dqm[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector151~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_3),
	.prn(vcc));
defparam \m_dqm[3] .is_wysiwyg = "true";
defparam \m_dqm[3] .power_up = "low";

dffeas \m_cmd[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_2),
	.prn(vcc));
defparam \m_cmd[2] .is_wysiwyg = "true";
defparam \m_cmd[2] .power_up = "low";

dffeas \m_cmd[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector22~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_0),
	.prn(vcc));
defparam \m_cmd[0] .is_wysiwyg = "true";
defparam \m_cmd[0] .power_up = "low";

dffeas \m_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector150~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_0),
	.prn(vcc));
defparam \m_data[0] .is_wysiwyg = "true";
defparam \m_data[0] .power_up = "low";

dffeas \m_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector149~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_1),
	.prn(vcc));
defparam \m_data[1] .is_wysiwyg = "true";
defparam \m_data[1] .power_up = "low";

dffeas \m_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector148~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_2),
	.prn(vcc));
defparam \m_data[2] .is_wysiwyg = "true";
defparam \m_data[2] .power_up = "low";

dffeas \m_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector147~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_3),
	.prn(vcc));
defparam \m_data[3] .is_wysiwyg = "true";
defparam \m_data[3] .power_up = "low";

dffeas \m_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\Selector146~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_4),
	.prn(vcc));
defparam \m_data[4] .is_wysiwyg = "true";
defparam \m_data[4] .power_up = "low";

dffeas \m_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\Selector145~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_5),
	.prn(vcc));
defparam \m_data[5] .is_wysiwyg = "true";
defparam \m_data[5] .power_up = "low";

dffeas \m_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\Selector144~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_6),
	.prn(vcc));
defparam \m_data[6] .is_wysiwyg = "true";
defparam \m_data[6] .power_up = "low";

dffeas \m_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\Selector143~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_7),
	.prn(vcc));
defparam \m_data[7] .is_wysiwyg = "true";
defparam \m_data[7] .power_up = "low";

dffeas \m_data[8] (
	.clk(wire_pll7_clk_0),
	.d(\Selector142~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_8),
	.prn(vcc));
defparam \m_data[8] .is_wysiwyg = "true";
defparam \m_data[8] .power_up = "low";

dffeas \m_data[9] (
	.clk(wire_pll7_clk_0),
	.d(\Selector141~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_9),
	.prn(vcc));
defparam \m_data[9] .is_wysiwyg = "true";
defparam \m_data[9] .power_up = "low";

dffeas \m_data[10] (
	.clk(wire_pll7_clk_0),
	.d(\Selector140~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_10),
	.prn(vcc));
defparam \m_data[10] .is_wysiwyg = "true";
defparam \m_data[10] .power_up = "low";

dffeas \m_data[11] (
	.clk(wire_pll7_clk_0),
	.d(\Selector139~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_11),
	.prn(vcc));
defparam \m_data[11] .is_wysiwyg = "true";
defparam \m_data[11] .power_up = "low";

dffeas \m_data[12] (
	.clk(wire_pll7_clk_0),
	.d(\Selector138~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_12),
	.prn(vcc));
defparam \m_data[12] .is_wysiwyg = "true";
defparam \m_data[12] .power_up = "low";

dffeas \m_data[13] (
	.clk(wire_pll7_clk_0),
	.d(\Selector137~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_13),
	.prn(vcc));
defparam \m_data[13] .is_wysiwyg = "true";
defparam \m_data[13] .power_up = "low";

dffeas \m_data[14] (
	.clk(wire_pll7_clk_0),
	.d(\Selector136~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_14),
	.prn(vcc));
defparam \m_data[14] .is_wysiwyg = "true";
defparam \m_data[14] .power_up = "low";

dffeas \m_data[15] (
	.clk(wire_pll7_clk_0),
	.d(\Selector135~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_15),
	.prn(vcc));
defparam \m_data[15] .is_wysiwyg = "true";
defparam \m_data[15] .power_up = "low";

dffeas \m_data[16] (
	.clk(wire_pll7_clk_0),
	.d(\Selector134~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_16),
	.prn(vcc));
defparam \m_data[16] .is_wysiwyg = "true";
defparam \m_data[16] .power_up = "low";

dffeas \m_data[17] (
	.clk(wire_pll7_clk_0),
	.d(\Selector133~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_17),
	.prn(vcc));
defparam \m_data[17] .is_wysiwyg = "true";
defparam \m_data[17] .power_up = "low";

dffeas \m_data[18] (
	.clk(wire_pll7_clk_0),
	.d(\Selector132~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_18),
	.prn(vcc));
defparam \m_data[18] .is_wysiwyg = "true";
defparam \m_data[18] .power_up = "low";

dffeas \m_data[19] (
	.clk(wire_pll7_clk_0),
	.d(\Selector131~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_19),
	.prn(vcc));
defparam \m_data[19] .is_wysiwyg = "true";
defparam \m_data[19] .power_up = "low";

dffeas \m_data[20] (
	.clk(wire_pll7_clk_0),
	.d(\Selector130~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_20),
	.prn(vcc));
defparam \m_data[20] .is_wysiwyg = "true";
defparam \m_data[20] .power_up = "low";

dffeas \m_data[21] (
	.clk(wire_pll7_clk_0),
	.d(\Selector129~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_21),
	.prn(vcc));
defparam \m_data[21] .is_wysiwyg = "true";
defparam \m_data[21] .power_up = "low";

dffeas \m_data[22] (
	.clk(wire_pll7_clk_0),
	.d(\Selector128~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_22),
	.prn(vcc));
defparam \m_data[22] .is_wysiwyg = "true";
defparam \m_data[22] .power_up = "low";

dffeas \m_data[23] (
	.clk(wire_pll7_clk_0),
	.d(\Selector127~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_23),
	.prn(vcc));
defparam \m_data[23] .is_wysiwyg = "true";
defparam \m_data[23] .power_up = "low";

dffeas \m_data[24] (
	.clk(wire_pll7_clk_0),
	.d(\Selector126~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_24),
	.prn(vcc));
defparam \m_data[24] .is_wysiwyg = "true";
defparam \m_data[24] .power_up = "low";

dffeas \m_data[25] (
	.clk(wire_pll7_clk_0),
	.d(\Selector125~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_25),
	.prn(vcc));
defparam \m_data[25] .is_wysiwyg = "true";
defparam \m_data[25] .power_up = "low";

dffeas \m_data[26] (
	.clk(wire_pll7_clk_0),
	.d(\Selector124~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_26),
	.prn(vcc));
defparam \m_data[26] .is_wysiwyg = "true";
defparam \m_data[26] .power_up = "low";

dffeas \m_data[27] (
	.clk(wire_pll7_clk_0),
	.d(\Selector123~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_27),
	.prn(vcc));
defparam \m_data[27] .is_wysiwyg = "true";
defparam \m_data[27] .power_up = "low";

dffeas \m_data[28] (
	.clk(wire_pll7_clk_0),
	.d(\Selector122~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_28),
	.prn(vcc));
defparam \m_data[28] .is_wysiwyg = "true";
defparam \m_data[28] .power_up = "low";

dffeas \m_data[29] (
	.clk(wire_pll7_clk_0),
	.d(\Selector121~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_29),
	.prn(vcc));
defparam \m_data[29] .is_wysiwyg = "true";
defparam \m_data[29] .power_up = "low";

dffeas \m_data[30] (
	.clk(wire_pll7_clk_0),
	.d(\Selector120~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_30),
	.prn(vcc));
defparam \m_data[30] .is_wysiwyg = "true";
defparam \m_data[30] .power_up = "low";

dffeas \m_data[31] (
	.clk(wire_pll7_clk_0),
	.d(\Selector119~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_31),
	.prn(vcc));
defparam \m_data[31] .is_wysiwyg = "true";
defparam \m_data[31] .power_up = "low";

dffeas za_valid(
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[2]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_valid1),
	.prn(vcc));
defparam za_valid.is_wysiwyg = "true";
defparam za_valid.power_up = "low";

dffeas \za_data[0] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_0),
	.prn(vcc));
defparam \za_data[0] .is_wysiwyg = "true";
defparam \za_data[0] .power_up = "low";

dffeas \za_data[1] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_1),
	.prn(vcc));
defparam \za_data[1] .is_wysiwyg = "true";
defparam \za_data[1] .power_up = "low";

dffeas \za_data[2] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_2),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_2),
	.prn(vcc));
defparam \za_data[2] .is_wysiwyg = "true";
defparam \za_data[2] .power_up = "low";

dffeas \za_data[3] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_3),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_3),
	.prn(vcc));
defparam \za_data[3] .is_wysiwyg = "true";
defparam \za_data[3] .power_up = "low";

dffeas \za_data[4] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_4),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_4),
	.prn(vcc));
defparam \za_data[4] .is_wysiwyg = "true";
defparam \za_data[4] .power_up = "low";

dffeas \za_data[22] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_22),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_22),
	.prn(vcc));
defparam \za_data[22] .is_wysiwyg = "true";
defparam \za_data[22] .power_up = "low";

dffeas \za_data[23] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_23),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_23),
	.prn(vcc));
defparam \za_data[23] .is_wysiwyg = "true";
defparam \za_data[23] .power_up = "low";

dffeas \za_data[24] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_24),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_24),
	.prn(vcc));
defparam \za_data[24] .is_wysiwyg = "true";
defparam \za_data[24] .power_up = "low";

dffeas \za_data[25] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_25),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_25),
	.prn(vcc));
defparam \za_data[25] .is_wysiwyg = "true";
defparam \za_data[25] .power_up = "low";

dffeas \za_data[26] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_26),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_26),
	.prn(vcc));
defparam \za_data[26] .is_wysiwyg = "true";
defparam \za_data[26] .power_up = "low";

dffeas \za_data[11] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_11),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_11),
	.prn(vcc));
defparam \za_data[11] .is_wysiwyg = "true";
defparam \za_data[11] .power_up = "low";

dffeas \za_data[13] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_13),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_13),
	.prn(vcc));
defparam \za_data[13] .is_wysiwyg = "true";
defparam \za_data[13] .power_up = "low";

dffeas \za_data[16] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_16),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_16),
	.prn(vcc));
defparam \za_data[16] .is_wysiwyg = "true";
defparam \za_data[16] .power_up = "low";

dffeas \za_data[12] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_12),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_12),
	.prn(vcc));
defparam \za_data[12] .is_wysiwyg = "true";
defparam \za_data[12] .power_up = "low";

dffeas \za_data[5] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_5),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_5),
	.prn(vcc));
defparam \za_data[5] .is_wysiwyg = "true";
defparam \za_data[5] .power_up = "low";

dffeas \za_data[14] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_14),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_14),
	.prn(vcc));
defparam \za_data[14] .is_wysiwyg = "true";
defparam \za_data[14] .power_up = "low";

dffeas \za_data[15] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_15),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_15),
	.prn(vcc));
defparam \za_data[15] .is_wysiwyg = "true";
defparam \za_data[15] .power_up = "low";

dffeas \za_data[10] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_10),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_10),
	.prn(vcc));
defparam \za_data[10] .is_wysiwyg = "true";
defparam \za_data[10] .power_up = "low";

dffeas \za_data[9] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_9),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_9),
	.prn(vcc));
defparam \za_data[9] .is_wysiwyg = "true";
defparam \za_data[9] .power_up = "low";

dffeas \za_data[8] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_8),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_8),
	.prn(vcc));
defparam \za_data[8] .is_wysiwyg = "true";
defparam \za_data[8] .power_up = "low";

dffeas \za_data[7] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_7),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_7),
	.prn(vcc));
defparam \za_data[7] .is_wysiwyg = "true";
defparam \za_data[7] .power_up = "low";

dffeas \za_data[6] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_6),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_6),
	.prn(vcc));
defparam \za_data[6] .is_wysiwyg = "true";
defparam \za_data[6] .power_up = "low";

dffeas \za_data[20] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_20),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_20),
	.prn(vcc));
defparam \za_data[20] .is_wysiwyg = "true";
defparam \za_data[20] .power_up = "low";

dffeas \za_data[18] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_18),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_18),
	.prn(vcc));
defparam \za_data[18] .is_wysiwyg = "true";
defparam \za_data[18] .power_up = "low";

dffeas \za_data[19] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_19),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_19),
	.prn(vcc));
defparam \za_data[19] .is_wysiwyg = "true";
defparam \za_data[19] .power_up = "low";

dffeas \za_data[17] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_17),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_17),
	.prn(vcc));
defparam \za_data[17] .is_wysiwyg = "true";
defparam \za_data[17] .power_up = "low";

dffeas \za_data[21] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_21),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_21),
	.prn(vcc));
defparam \za_data[21] .is_wysiwyg = "true";
defparam \za_data[21] .power_up = "low";

dffeas \za_data[27] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_27),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_27),
	.prn(vcc));
defparam \za_data[27] .is_wysiwyg = "true";
defparam \za_data[27] .power_up = "low";

dffeas \za_data[28] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_28),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_28),
	.prn(vcc));
defparam \za_data[28] .is_wysiwyg = "true";
defparam \za_data[28] .power_up = "low";

dffeas \za_data[31] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_31),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_31),
	.prn(vcc));
defparam \za_data[31] .is_wysiwyg = "true";
defparam \za_data[31] .power_up = "low";

dffeas \za_data[30] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_30),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_30),
	.prn(vcc));
defparam \za_data[30] .is_wysiwyg = "true";
defparam \za_data[30] .power_up = "low";

dffeas \za_data[29] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_29),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_29),
	.prn(vcc));
defparam \za_data[29] .is_wysiwyg = "true";
defparam \za_data[29] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\refresh_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh_counter~9 (
	.dataa(\Add0~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~9_combout ),
	.cout());
defparam \refresh_counter~9 .lut_mask = 16'hAAFF;
defparam \refresh_counter~9 .sum_lutc_input = "datac";

dffeas \refresh_counter[0] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[0]~q ),
	.prn(vcc));
defparam \refresh_counter[0] .is_wysiwyg = "true";
defparam \refresh_counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\refresh_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

dffeas \refresh_counter[1] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[1]~q ),
	.prn(vcc));
defparam \refresh_counter[1] .is_wysiwyg = "true";
defparam \refresh_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add0~4 (
	.dataa(\refresh_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

dffeas \refresh_counter[2] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[2]~q ),
	.prn(vcc));
defparam \refresh_counter[2] .is_wysiwyg = "true";
defparam \refresh_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add0~6 (
	.dataa(\refresh_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~8 (
	.dataa(\Add0~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~8_combout ),
	.cout());
defparam \refresh_counter~8 .lut_mask = 16'hAAFF;
defparam \refresh_counter~8 .sum_lutc_input = "datac";

dffeas \refresh_counter[3] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[3]~q ),
	.prn(vcc));
defparam \refresh_counter[3] .is_wysiwyg = "true";
defparam \refresh_counter[3] .power_up = "low";

cycloneive_lcell_comb \Add0~8 (
	.dataa(\refresh_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~6 (
	.dataa(\Add0~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~6_combout ),
	.cout());
defparam \refresh_counter~6 .lut_mask = 16'hFF55;
defparam \refresh_counter~6 .sum_lutc_input = "datac";

dffeas \refresh_counter[4] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[4]~q ),
	.prn(vcc));
defparam \refresh_counter[4] .is_wysiwyg = "true";
defparam \refresh_counter[4] .power_up = "low";

cycloneive_lcell_comb \Add0~10 (
	.dataa(\refresh_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~7 (
	.dataa(\Add0~10_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~7_combout ),
	.cout());
defparam \refresh_counter~7 .lut_mask = 16'hAAFF;
defparam \refresh_counter~7 .sum_lutc_input = "datac";

dffeas \refresh_counter[5] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[5]~q ),
	.prn(vcc));
defparam \refresh_counter[5] .is_wysiwyg = "true";
defparam \refresh_counter[5] .power_up = "low";

cycloneive_lcell_comb \Add0~12 (
	.dataa(\refresh_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~5 (
	.dataa(\Add0~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~5_combout ),
	.cout());
defparam \refresh_counter~5 .lut_mask = 16'hAAFF;
defparam \refresh_counter~5 .sum_lutc_input = "datac";

dffeas \refresh_counter[6] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[6]~q ),
	.prn(vcc));
defparam \refresh_counter[6] .is_wysiwyg = "true";
defparam \refresh_counter[6] .power_up = "low";

cycloneive_lcell_comb \Add0~14 (
	.dataa(\refresh_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

dffeas \refresh_counter[7] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~14_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[7]~q ),
	.prn(vcc));
defparam \refresh_counter[7] .is_wysiwyg = "true";
defparam \refresh_counter[7] .power_up = "low";

cycloneive_lcell_comb \Add0~16 (
	.dataa(\refresh_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'h5A5F;
defparam \Add0~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter[8]~13 (
	.dataa(\Add0~16_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\refresh_counter[8]~13_combout ),
	.cout());
defparam \refresh_counter[8]~13 .lut_mask = 16'h5555;
defparam \refresh_counter[8]~13 .sum_lutc_input = "datac";

dffeas \refresh_counter[8] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter[8]~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[8]~q ),
	.prn(vcc));
defparam \refresh_counter[8] .is_wysiwyg = "true";
defparam \refresh_counter[8] .power_up = "low";

cycloneive_lcell_comb \Add0~18 (
	.dataa(\refresh_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'h5AAF;
defparam \Add0~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~4 (
	.dataa(\Add0~18_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~4_combout ),
	.cout());
defparam \refresh_counter~4 .lut_mask = 16'hFF55;
defparam \refresh_counter~4 .sum_lutc_input = "datac";

dffeas \refresh_counter[9] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[9]~q ),
	.prn(vcc));
defparam \refresh_counter[9] .is_wysiwyg = "true";
defparam \refresh_counter[9] .power_up = "low";

cycloneive_lcell_comb \Add0~20 (
	.dataa(\refresh_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h5A5F;
defparam \Add0~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~1 (
	.dataa(\Add0~20_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~1_combout ),
	.cout());
defparam \refresh_counter~1 .lut_mask = 16'hFF55;
defparam \refresh_counter~1 .sum_lutc_input = "datac";

dffeas \refresh_counter[10] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[10]~q ),
	.prn(vcc));
defparam \refresh_counter[10] .is_wysiwyg = "true";
defparam \refresh_counter[10] .power_up = "low";

cycloneive_lcell_comb \Add0~22 (
	.dataa(\refresh_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~3 (
	.dataa(\Add0~22_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~3_combout ),
	.cout());
defparam \refresh_counter~3 .lut_mask = 16'hAAFF;
defparam \refresh_counter~3 .sum_lutc_input = "datac";

dffeas \refresh_counter[11] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[11]~q ),
	.prn(vcc));
defparam \refresh_counter[11] .is_wysiwyg = "true";
defparam \refresh_counter[11] .power_up = "low";

cycloneive_lcell_comb \Add0~24 (
	.dataa(\refresh_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'h5AAF;
defparam \Add0~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~2 (
	.dataa(\Add0~24_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~2_combout ),
	.cout());
defparam \refresh_counter~2 .lut_mask = 16'hAAFF;
defparam \refresh_counter~2 .sum_lutc_input = "datac";

dffeas \refresh_counter[12] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[12]~q ),
	.prn(vcc));
defparam \refresh_counter[12] .is_wysiwyg = "true";
defparam \refresh_counter[12] .power_up = "low";

cycloneive_lcell_comb \Add0~26 (
	.dataa(\refresh_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout());
defparam \Add0~26 .lut_mask = 16'h5A5A;
defparam \Add0~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~0 (
	.dataa(\Add0~26_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~0_combout ),
	.cout());
defparam \refresh_counter~0 .lut_mask = 16'hFF55;
defparam \refresh_counter~0 .sum_lutc_input = "datac";

dffeas \refresh_counter[13] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[13]~q ),
	.prn(vcc));
defparam \refresh_counter[13] .is_wysiwyg = "true";
defparam \refresh_counter[13] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\refresh_counter[13]~q ),
	.datab(\refresh_counter[10]~q ),
	.datac(\refresh_counter[12]~q ),
	.datad(\refresh_counter[11]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\refresh_counter[9]~q ),
	.datab(\refresh_counter[8]~q ),
	.datac(\refresh_counter[7]~q ),
	.datad(\refresh_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\refresh_counter[4]~q ),
	.datab(\refresh_counter[5]~q ),
	.datac(\refresh_counter[3]~q ),
	.datad(\refresh_counter[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hBFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\refresh_counter[1]~q ),
	.datad(\refresh_counter[0]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h0FFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hFFFE;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_next.000~0 (
	.dataa(\i_next.000~q ),
	.datab(\i_state.000~q ),
	.datac(\i_state.101~q ),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\i_next.000~0_combout ),
	.cout());
defparam \i_next.000~0 .lut_mask = 16'hEFFF;
defparam \i_next.000~0 .sum_lutc_input = "datac";

dffeas \i_next.000 (
	.clk(wire_pll7_clk_0),
	.d(\i_next.000~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.000~q ),
	.prn(vcc));
defparam \i_next.000 .is_wysiwyg = "true";
defparam \i_next.000 .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\i_count[0]~0_combout ),
	.datab(\i_state.000~q ),
	.datac(\Equal0~4_combout ),
	.datad(\i_next.000~q ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFFFD;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \i_state.000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.000~q ),
	.prn(vcc));
defparam \i_state.000 .is_wysiwyg = "true";
defparam \i_state.000 .power_up = "low";

cycloneive_lcell_comb \Selector18~0 (
	.dataa(\i_next.111~q ),
	.datab(\i_state.101~q ),
	.datac(\i_state.011~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
defparam \Selector18~0 .lut_mask = 16'hFEFF;
defparam \Selector18~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hAAFF;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \i_state.001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.001~q ),
	.prn(vcc));
defparam \i_state.001 .is_wysiwyg = "true";
defparam \i_state.001 .power_up = "low";

cycloneive_lcell_comb \Selector16~0 (
	.dataa(\i_next.010~q ),
	.datab(\i_state.101~q ),
	.datac(\i_state.011~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
defparam \Selector16~0 .lut_mask = 16'hFEFF;
defparam \Selector16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(\i_state.010~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hAFFA;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas \i_refs[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(altera_reset_synchronizer_int_chain_out),
	.q(\i_refs[0]~q ),
	.prn(vcc));
defparam \i_refs[0] .is_wysiwyg = "true";
defparam \i_refs[0] .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\i_state.000~q ),
	.datab(\i_state.010~q ),
	.datac(\i_refs[1]~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEBBE;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \i_refs[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(altera_reset_synchronizer_int_chain_out),
	.q(\i_refs[1]~q ),
	.prn(vcc));
defparam \i_refs[1] .is_wysiwyg = "true";
defparam \i_refs[1] .power_up = "low";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\i_state.010~q ),
	.datab(\i_refs[2]~q ),
	.datac(\i_refs[1]~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEBBE;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(\Selector4~0_combout ),
	.datab(\i_state.000~q ),
	.datac(\i_refs[2]~q ),
	.datad(\i_state.010~q ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hFEFF;
defparam \Selector4~1 .sum_lutc_input = "datac";

dffeas \i_refs[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(altera_reset_synchronizer_int_chain_out),
	.q(\i_refs[2]~q ),
	.prn(vcc));
defparam \i_refs[2] .is_wysiwyg = "true";
defparam \i_refs[2] .power_up = "low";

cycloneive_lcell_comb \Selector18~1 (
	.dataa(\i_refs[0]~q ),
	.datab(gnd),
	.datac(\i_refs[2]~q ),
	.datad(\i_refs[1]~q ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
defparam \Selector18~1 .lut_mask = 16'hAFFF;
defparam \Selector18~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector16~1 (
	.dataa(\i_state.001~q ),
	.datab(\Selector16~0_combout ),
	.datac(\i_state.010~q ),
	.datad(\Selector18~1_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
defparam \Selector16~1 .lut_mask = 16'hFEFF;
defparam \Selector16~1 .sum_lutc_input = "datac";

dffeas \i_next.010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector16~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.010~q ),
	.prn(vcc));
defparam \i_next.010 .is_wysiwyg = "true";
defparam \i_next.010 .power_up = "low";

cycloneive_lcell_comb \i_count[0]~4 (
	.dataa(\i_state.010~q ),
	.datab(gnd),
	.datac(\i_state.011~q ),
	.datad(\i_count[0]~q ),
	.cin(gnd),
	.combout(\i_count[0]~4_combout ),
	.cout());
defparam \i_count[0]~4 .lut_mask = 16'hA0AF;
defparam \i_count[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_count[0]~1 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.101~q ),
	.cin(gnd),
	.combout(\i_count[0]~1_combout ),
	.cout());
defparam \i_count[0]~1 .lut_mask = 16'hAAFF;
defparam \i_count[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_count[0]~5 (
	.dataa(\i_count[0]~q ),
	.datab(\i_count[0]~4_combout ),
	.datac(\i_count[0]~1_combout ),
	.datad(\i_count[0]~0_combout ),
	.cin(gnd),
	.combout(\i_count[0]~5_combout ),
	.cout());
defparam \i_count[0]~5 .lut_mask = 16'hEFFE;
defparam \i_count[0]~5 .sum_lutc_input = "datac";

dffeas \i_count[0] (
	.clk(wire_pll7_clk_0),
	.d(\i_count[0]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[0]~q ),
	.prn(vcc));
defparam \i_count[0] .is_wysiwyg = "true";
defparam \i_count[0] .power_up = "low";

cycloneive_lcell_comb \i_count[1]~2 (
	.dataa(\i_count[1]~q ),
	.datab(\i_count[0]~q ),
	.datac(\i_state.010~q ),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\i_count[1]~2_combout ),
	.cout());
defparam \i_count[1]~2 .lut_mask = 16'hF9F6;
defparam \i_count[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_count[1]~3 (
	.dataa(\i_count[1]~q ),
	.datab(\i_count[1]~2_combout ),
	.datac(\i_count[0]~1_combout ),
	.datad(\i_count[0]~0_combout ),
	.cin(gnd),
	.combout(\i_count[1]~3_combout ),
	.cout());
defparam \i_count[1]~3 .lut_mask = 16'hEFFE;
defparam \i_count[1]~3 .sum_lutc_input = "datac";

dffeas \i_count[1] (
	.clk(wire_pll7_clk_0),
	.d(\i_count[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[1]~q ),
	.prn(vcc));
defparam \i_count[1] .is_wysiwyg = "true";
defparam \i_count[1] .power_up = "low";

cycloneive_lcell_comb \Selector13~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_count[1]~q ),
	.datac(\i_count[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hFEFE;
defparam \Selector13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector13~1 (
	.dataa(\i_state.111~q ),
	.datab(\i_count[2]~q ),
	.datac(\Selector13~0_combout ),
	.datad(\i_count[0]~1_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
defparam \Selector13~1 .lut_mask = 16'hFEFF;
defparam \Selector13~1 .sum_lutc_input = "datac";

dffeas \i_count[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector13~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[2]~q ),
	.prn(vcc));
defparam \i_count[2] .is_wysiwyg = "true";
defparam \i_count[2] .power_up = "low";

cycloneive_lcell_comb \Selector9~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_next.010~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hEFFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

dffeas \i_state.010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.010~q ),
	.prn(vcc));
defparam \i_state.010 .is_wysiwyg = "true";
defparam \i_state.010 .power_up = "low";

cycloneive_lcell_comb \Selector18~2 (
	.dataa(\Selector18~0_combout ),
	.datab(\i_state.010~q ),
	.datac(\Selector18~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
defparam \Selector18~2 .lut_mask = 16'hFEFE;
defparam \Selector18~2 .sum_lutc_input = "datac";

dffeas \i_next.111 (
	.clk(wire_pll7_clk_0),
	.d(\Selector18~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.111~q ),
	.prn(vcc));
defparam \i_next.111 .is_wysiwyg = "true";
defparam \i_next.111 .power_up = "low";

cycloneive_lcell_comb \Selector12~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_next.111~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'hEFFF;
defparam \Selector12~0 .sum_lutc_input = "datac";

dffeas \i_state.111 (
	.clk(wire_pll7_clk_0),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.111~q ),
	.prn(vcc));
defparam \i_state.111 .is_wysiwyg = "true";
defparam \i_state.111 .power_up = "low";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(\i_state.001~q ),
	.datab(\i_state.011~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFFFE;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~1 (
	.dataa(\i_state.111~q ),
	.datab(\i_state.010~q ),
	.datac(\Selector10~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hFEFE;
defparam \Selector10~1 .sum_lutc_input = "datac";

dffeas \i_state.011 (
	.clk(wire_pll7_clk_0),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.011~q ),
	.prn(vcc));
defparam \i_state.011 .is_wysiwyg = "true";
defparam \i_state.011 .power_up = "low";

cycloneive_lcell_comb \i_count[0]~0 (
	.dataa(\i_state.011~q ),
	.datab(gnd),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\i_count[0]~0_combout ),
	.cout());
defparam \i_count[0]~0 .lut_mask = 16'hAFFF;
defparam \i_count[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr6~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\WideOr6~0_combout ),
	.cout());
defparam \WideOr6~0 .lut_mask = 16'hAAFF;
defparam \WideOr6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector17~0 (
	.dataa(\i_state.111~q ),
	.datab(\i_next.101~q ),
	.datac(\i_state.101~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
defparam \Selector17~0 .lut_mask = 16'hFEFF;
defparam \Selector17~0 .sum_lutc_input = "datac";

dffeas \i_next.101 (
	.clk(wire_pll7_clk_0),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.101~q ),
	.prn(vcc));
defparam \i_next.101 .is_wysiwyg = "true";
defparam \i_next.101 .power_up = "low";

cycloneive_lcell_comb \i_state.101~0 (
	.dataa(\i_state.101~q ),
	.datab(\i_count[0]~0_combout ),
	.datac(\i_next.101~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\i_state.101~0_combout ),
	.cout());
defparam \i_state.101~0 .lut_mask = 16'hFEFE;
defparam \i_state.101~0 .sum_lutc_input = "datac";

dffeas \i_state.101 (
	.clk(wire_pll7_clk_0),
	.d(\i_state.101~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.101~q ),
	.prn(vcc));
defparam \i_state.101 .is_wysiwyg = "true";
defparam \i_state.101 .power_up = "low";

cycloneive_lcell_comb \init_done~0 (
	.dataa(\init_done~q ),
	.datab(\i_state.101~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\init_done~0_combout ),
	.cout());
defparam \init_done~0 .lut_mask = 16'hEEEE;
defparam \init_done~0 .sum_lutc_input = "datac";

dffeas init_done(
	.clk(wire_pll7_clk_0),
	.d(\init_done~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\init_done~q ),
	.prn(vcc));
defparam init_done.is_wysiwyg = "true";
defparam init_done.power_up = "low";

cycloneive_lcell_comb \Selector24~1 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\refresh_request~q ),
	.datad(\init_done~q ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
defparam \Selector24~1 .lut_mask = 16'h7FFF;
defparam \Selector24~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~0 (
	.dataa(\m_state.100000000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector32~0_combout ),
	.cout());
defparam \Selector32~0 .lut_mask = 16'hAAFF;
defparam \Selector32~0 .sum_lutc_input = "datac";

dffeas active_rnw(
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_rnw~q ),
	.prn(vcc));
defparam active_rnw.is_wysiwyg = "true";
defparam active_rnw.power_up = "low";

cycloneive_lcell_comb \Selector25~5 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(gnd),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
defparam \Selector25~5 .lut_mask = 16'hEEFF;
defparam \Selector25~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector25~6 (
	.dataa(\init_done~q ),
	.datab(\m_state.000000001~q ),
	.datac(\Selector25~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector25~6_combout ),
	.cout());
defparam \Selector25~6 .lut_mask = 16'hFBFB;
defparam \Selector25~6 .sum_lutc_input = "datac";

dffeas \m_state.000000010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector25~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000010~q ),
	.prn(vcc));
defparam \m_state.000000010 .is_wysiwyg = "true";
defparam \m_state.000000010 .power_up = "low";

dffeas \active_addr[10] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[10]~q ),
	.prn(vcc));
defparam \active_addr[10] .is_wysiwyg = "true";
defparam \active_addr[10] .power_up = "low";

cycloneive_lcell_comb \pending~0 (
	.dataa(\active_rnw~q ),
	.datab(\active_addr[10]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.cin(gnd),
	.combout(\pending~0_combout ),
	.cout());
defparam \pending~0 .lut_mask = 16'h6996;
defparam \pending~0 .sum_lutc_input = "datac";

dffeas \active_addr[24] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[24]~q ),
	.prn(vcc));
defparam \active_addr[24] .is_wysiwyg = "true";
defparam \active_addr[24] .power_up = "low";

cycloneive_lcell_comb \pending~1 (
	.dataa(\active_addr[11]~q ),
	.datab(\active_addr[24]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[47]~3_combout ),
	.cin(gnd),
	.combout(\pending~1_combout ),
	.cout());
defparam \pending~1 .lut_mask = 16'h6996;
defparam \pending~1 .sum_lutc_input = "datac";

dffeas \active_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[48]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[12]~q ),
	.prn(vcc));
defparam \active_addr[12] .is_wysiwyg = "true";
defparam \active_addr[12] .power_up = "low";

dffeas \active_addr[13] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[49]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[13]~q ),
	.prn(vcc));
defparam \active_addr[13] .is_wysiwyg = "true";
defparam \active_addr[13] .power_up = "low";

cycloneive_lcell_comb \pending~2 (
	.dataa(\active_addr[12]~q ),
	.datab(\active_addr[13]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[49]~4_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[48]~5_combout ),
	.cin(gnd),
	.combout(\pending~2_combout ),
	.cout());
defparam \pending~2 .lut_mask = 16'h6996;
defparam \pending~2 .sum_lutc_input = "datac";

dffeas \active_addr[14] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[50]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[14]~q ),
	.prn(vcc));
defparam \active_addr[14] .is_wysiwyg = "true";
defparam \active_addr[14] .power_up = "low";

dffeas \active_addr[15] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[51]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[15]~q ),
	.prn(vcc));
defparam \active_addr[15] .is_wysiwyg = "true";
defparam \active_addr[15] .power_up = "low";

cycloneive_lcell_comb \pending~3 (
	.dataa(\active_addr[14]~q ),
	.datab(\active_addr[15]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[51]~6_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[50]~7_combout ),
	.cin(gnd),
	.combout(\pending~3_combout ),
	.cout());
defparam \pending~3 .lut_mask = 16'h6996;
defparam \pending~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~4 (
	.dataa(\pending~0_combout ),
	.datab(\pending~1_combout ),
	.datac(\pending~2_combout ),
	.datad(\pending~3_combout ),
	.cin(gnd),
	.combout(\pending~4_combout ),
	.cout());
defparam \pending~4 .lut_mask = 16'hFFFE;
defparam \pending~4 .sum_lutc_input = "datac";

dffeas \active_addr[16] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[52]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[16]~q ),
	.prn(vcc));
defparam \active_addr[16] .is_wysiwyg = "true";
defparam \active_addr[16] .power_up = "low";

dffeas \active_addr[17] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[53]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[17]~q ),
	.prn(vcc));
defparam \active_addr[17] .is_wysiwyg = "true";
defparam \active_addr[17] .power_up = "low";

cycloneive_lcell_comb \pending~5 (
	.dataa(\active_addr[16]~q ),
	.datab(\active_addr[17]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[53]~8_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[52]~9_combout ),
	.cin(gnd),
	.combout(\pending~5_combout ),
	.cout());
defparam \pending~5 .lut_mask = 16'h6996;
defparam \pending~5 .sum_lutc_input = "datac";

dffeas \active_addr[18] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[54]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[18]~q ),
	.prn(vcc));
defparam \active_addr[18] .is_wysiwyg = "true";
defparam \active_addr[18] .power_up = "low";

dffeas \active_addr[19] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[55]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[19]~q ),
	.prn(vcc));
defparam \active_addr[19] .is_wysiwyg = "true";
defparam \active_addr[19] .power_up = "low";

cycloneive_lcell_comb \pending~6 (
	.dataa(\active_addr[18]~q ),
	.datab(\active_addr[19]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[55]~10_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[54]~11_combout ),
	.cin(gnd),
	.combout(\pending~6_combout ),
	.cout());
defparam \pending~6 .lut_mask = 16'h6996;
defparam \pending~6 .sum_lutc_input = "datac";

dffeas \active_addr[20] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[56]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[20]~q ),
	.prn(vcc));
defparam \active_addr[20] .is_wysiwyg = "true";
defparam \active_addr[20] .power_up = "low";

dffeas \active_addr[21] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[57]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[21]~q ),
	.prn(vcc));
defparam \active_addr[21] .is_wysiwyg = "true";
defparam \active_addr[21] .power_up = "low";

cycloneive_lcell_comb \pending~7 (
	.dataa(\active_addr[20]~q ),
	.datab(\active_addr[21]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[57]~12_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[56]~13_combout ),
	.cin(gnd),
	.combout(\pending~7_combout ),
	.cout());
defparam \pending~7 .lut_mask = 16'h6996;
defparam \pending~7 .sum_lutc_input = "datac";

dffeas \active_addr[22] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[58]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[22]~q ),
	.prn(vcc));
defparam \active_addr[22] .is_wysiwyg = "true";
defparam \active_addr[22] .power_up = "low";

dffeas \active_addr[23] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[59]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[23]~q ),
	.prn(vcc));
defparam \active_addr[23] .is_wysiwyg = "true";
defparam \active_addr[23] .power_up = "low";

cycloneive_lcell_comb \pending~8 (
	.dataa(\active_addr[22]~q ),
	.datab(\active_addr[23]~q ),
	.datac(\the_usb_system_sdram_input_efifo_module|rd_data[59]~14_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[58]~15_combout ),
	.cin(gnd),
	.combout(\pending~8_combout ),
	.cout());
defparam \pending~8 .lut_mask = 16'h6996;
defparam \pending~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~9 (
	.dataa(\pending~5_combout ),
	.datab(\pending~6_combout ),
	.datac(\pending~7_combout ),
	.datad(\pending~8_combout ),
	.cin(gnd),
	.combout(\pending~9_combout ),
	.cout());
defparam \pending~9 .lut_mask = 16'hFFFE;
defparam \pending~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~10 (
	.dataa(\pending~4_combout ),
	.datab(\pending~9_combout ),
	.datac(gnd),
	.datad(\active_cs_n~q ),
	.cin(gnd),
	.combout(\pending~10_combout ),
	.cout());
defparam \pending~10 .lut_mask = 16'hEEFF;
defparam \pending~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_next~22 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\refresh_request~q ),
	.datad(\pending~10_combout ),
	.cin(gnd),
	.combout(\m_next~22_combout ),
	.cout());
defparam \m_next~22 .lut_mask = 16'hFEFF;
defparam \m_next~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector25~4 (
	.dataa(\init_done~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
defparam \Selector25~4 .lut_mask = 16'hAAFF;
defparam \Selector25~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~0 (
	.dataa(\m_state.100000000~q ),
	.datab(\pending~10_combout ),
	.datac(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hEFFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_next~21 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\pending~10_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\m_next~21_combout ),
	.cout());
defparam \m_next~21 .lut_mask = 16'hFFFE;
defparam \m_next~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector29~0 (
	.dataa(\m_state.100000000~q ),
	.datab(\active_cs_n~q ),
	.datac(\pending~4_combout ),
	.datad(\pending~9_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
defparam \Selector29~0 .lut_mask = 16'hEFFF;
defparam \Selector29~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~1 (
	.dataa(\m_count[0]~q ),
	.datab(\m_state.000000001~q ),
	.datac(\init_done~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector39~1_combout ),
	.cout());
defparam \Selector39~1 .lut_mask = 16'hEFFF;
defparam \Selector39~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~2 (
	.dataa(gnd),
	.datab(\m_state.000000100~q ),
	.datac(\m_count[1]~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector39~2_combout ),
	.cout());
defparam \Selector39~2 .lut_mask = 16'h3FFF;
defparam \Selector39~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~3 (
	.dataa(\Selector39~1_combout ),
	.datab(\Selector39~2_combout ),
	.datac(\m_state.000001000~q ),
	.datad(\m_next~21_combout ),
	.cin(gnd),
	.combout(\Selector39~3_combout ),
	.cout());
defparam \Selector39~3 .lut_mask = 16'hEFFF;
defparam \Selector39~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr10~0 (
	.dataa(\m_state.000000001~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_state.001000000~q ),
	.cin(gnd),
	.combout(\WideOr10~0_combout ),
	.cout());
defparam \WideOr10~0 .lut_mask = 16'hAAFF;
defparam \WideOr10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~0 (
	.dataa(\Selector24~0_combout ),
	.datab(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\refresh_request~q ),
	.datad(\m_state.100000000~q ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
defparam \Selector27~0 .lut_mask = 16'hBFFF;
defparam \Selector27~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~5 (
	.dataa(\Selector35~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\active_rnw~q ),
	.cin(gnd),
	.combout(\Selector35~5_combout ),
	.cout());
defparam \Selector35~5 .lut_mask = 16'hAAFF;
defparam \Selector35~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~1 (
	.dataa(\m_state.000000010~q ),
	.datab(\refresh_request~q ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector34~1_combout ),
	.cout());
defparam \Selector34~1 .lut_mask = 16'hEFFF;
defparam \Selector34~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~3 (
	.dataa(\m_state.100000000~q ),
	.datab(\m_state.010000000~q ),
	.datac(\refresh_request~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector35~3_combout ),
	.cout());
defparam \Selector35~3 .lut_mask = 16'h7F7F;
defparam \Selector35~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~4 (
	.dataa(\m_state.100000000~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\pending~10_combout ),
	.datad(\Selector35~3_combout ),
	.cin(gnd),
	.combout(\Selector35~4_combout ),
	.cout());
defparam \Selector35~4 .lut_mask = 16'hFFF7;
defparam \Selector35~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~2 (
	.dataa(\Selector34~1_combout ),
	.datab(\m_next~21_combout ),
	.datac(\WideOr9~0_combout ),
	.datad(\Selector35~4_combout ),
	.cin(gnd),
	.combout(\Selector34~2_combout ),
	.cout());
defparam \Selector34~2 .lut_mask = 16'hEFFF;
defparam \Selector34~2 .sum_lutc_input = "datac";

dffeas \m_next.000010000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector35~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector34~2_combout ),
	.q(\m_next.000010000~q ),
	.prn(vcc));
defparam \m_next.000010000 .is_wysiwyg = "true";
defparam \m_next.000010000 .power_up = "low";

cycloneive_lcell_comb \Selector27~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\pending~10_combout ),
	.datac(\m_state.100000000~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
defparam \Selector27~1 .lut_mask = 16'hFEFF;
defparam \Selector27~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector28~0 (
	.dataa(\Selector27~0_combout ),
	.datab(\m_next.000010000~q ),
	.datac(\Selector27~1_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
defparam \Selector28~0 .lut_mask = 16'hFEFF;
defparam \Selector28~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~3 (
	.dataa(\refresh_request~q ),
	.datab(\pending~combout ),
	.datac(\m_state.000000001~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
defparam \Selector27~3 .lut_mask = 16'hFEFF;
defparam \Selector27~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~4 (
	.dataa(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\refresh_request~q ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
defparam \Selector27~4 .lut_mask = 16'hEFFF;
defparam \Selector27~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr8~0 (
	.dataa(gnd),
	.datab(\m_state.000000010~q ),
	.datac(\m_state.001000000~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\WideOr8~0_combout ),
	.cout());
defparam \WideOr8~0 .lut_mask = 16'h3FFF;
defparam \WideOr8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~5 (
	.dataa(\m_state.100000000~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\refresh_request~q ),
	.datad(\WideOr8~0_combout ),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
defparam \Selector27~5 .lut_mask = 16'hFEFF;
defparam \Selector27~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~6 (
	.dataa(\Selector24~0_combout ),
	.datab(\Selector27~3_combout ),
	.datac(\Selector27~4_combout ),
	.datad(\Selector27~5_combout ),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
defparam \Selector27~6 .lut_mask = 16'hFFFE;
defparam \Selector27~6 .sum_lutc_input = "datac";

dffeas \m_state.000010000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector27~6_combout ),
	.q(\m_state.000010000~q ),
	.prn(vcc));
defparam \m_state.000010000 .is_wysiwyg = "true";
defparam \m_state.000010000 .power_up = "low";

cycloneive_lcell_comb \Selector39~0 (
	.dataa(\m_next~21_combout ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000001000~q ),
	.datad(\Selector38~0_combout ),
	.cin(gnd),
	.combout(\Selector39~0_combout ),
	.cout());
defparam \Selector39~0 .lut_mask = 16'hBFFF;
defparam \Selector39~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~4 (
	.dataa(\m_count[1]~q ),
	.datab(\m_state.000000100~q ),
	.datac(\m_state.000100000~q ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector39~4_combout ),
	.cout());
defparam \Selector39~4 .lut_mask = 16'hBFFF;
defparam \Selector39~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~5 (
	.dataa(\Selector39~3_combout ),
	.datab(\WideOr10~0_combout ),
	.datac(\Selector39~0_combout ),
	.datad(\Selector39~4_combout ),
	.cin(gnd),
	.combout(\Selector39~5_combout ),
	.cout());
defparam \Selector39~5 .lut_mask = 16'hFFFE;
defparam \Selector39~5 .sum_lutc_input = "datac";

dffeas \m_count[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector39~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[0]~q ),
	.prn(vcc));
defparam \m_count[0] .is_wysiwyg = "true";
defparam \m_count[0] .power_up = "low";

cycloneive_lcell_comb \Selector38~1 (
	.dataa(\m_count[1]~q ),
	.datab(\m_count[0]~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector38~1_combout ),
	.cout());
defparam \Selector38~1 .lut_mask = 16'hFFFE;
defparam \Selector38~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~2 (
	.dataa(\m_state.010000000~q ),
	.datab(\Selector38~1_combout ),
	.datac(\m_state.000001000~q ),
	.datad(\m_next~21_combout ),
	.cin(gnd),
	.combout(\Selector38~2_combout ),
	.cout());
defparam \Selector38~2 .lut_mask = 16'hFFFE;
defparam \Selector38~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~3 (
	.dataa(\m_state.001000000~q ),
	.datab(\init_done~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector38~3_combout ),
	.cout());
defparam \Selector38~3 .lut_mask = 16'hBFFF;
defparam \Selector38~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~4 (
	.dataa(\Selector38~2_combout ),
	.datab(\m_count[1]~q ),
	.datac(\Selector38~3_combout ),
	.datad(\Selector39~0_combout ),
	.cin(gnd),
	.combout(\Selector38~4_combout ),
	.cout());
defparam \Selector38~4 .lut_mask = 16'hFEFF;
defparam \Selector38~4 .sum_lutc_input = "datac";

dffeas \m_count[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector38~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[1]~q ),
	.prn(vcc));
defparam \m_count[1] .is_wysiwyg = "true";
defparam \m_count[1] .power_up = "low";

cycloneive_lcell_comb \Selector29~1 (
	.dataa(\m_state.000100000~q ),
	.datab(\Selector29~0_combout ),
	.datac(\Selector25~5_combout ),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
defparam \Selector29~1 .lut_mask = 16'hFFFE;
defparam \Selector29~1 .sum_lutc_input = "datac";

dffeas \m_state.000100000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector29~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000100000~q ),
	.prn(vcc));
defparam \m_state.000100000 .is_wysiwyg = "true";
defparam \m_state.000100000 .power_up = "low";

cycloneive_lcell_comb \Selector30~0 (
	.dataa(\m_state.000100000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
defparam \Selector30~0 .lut_mask = 16'hAAFF;
defparam \Selector30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector30~1 (
	.dataa(\Selector30~0_combout ),
	.datab(\init_done~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector30~1_combout ),
	.cout());
defparam \Selector30~1 .lut_mask = 16'hFEFF;
defparam \Selector30~1 .sum_lutc_input = "datac";

dffeas \m_state.001000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector30~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.001000000~q ),
	.prn(vcc));
defparam \m_state.001000000 .is_wysiwyg = "true";
defparam \m_state.001000000 .power_up = "low";

cycloneive_lcell_comb \Selector33~0 (
	.dataa(gnd),
	.datab(\m_state.001000000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector33~0_combout ),
	.cout());
defparam \Selector33~0 .lut_mask = 16'h3FFF;
defparam \Selector33~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~0 (
	.dataa(\Selector38~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\m_next~21_combout ),
	.datad(\Selector33~0_combout ),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
defparam \Selector36~0 .lut_mask = 16'hBFFF;
defparam \Selector36~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~1 (
	.dataa(\Selector25~4_combout ),
	.datab(\m_next.010000000~q ),
	.datac(\Selector36~0_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector36~1_combout ),
	.cout());
defparam \Selector36~1 .lut_mask = 16'hFFFE;
defparam \Selector36~1 .sum_lutc_input = "datac";

dffeas \m_next.010000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector36~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.010000000~q ),
	.prn(vcc));
defparam \m_next.010000000 .is_wysiwyg = "true";
defparam \m_next.010000000 .power_up = "low";

cycloneive_lcell_comb \Selector31~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_next.010000000~q ),
	.datac(gnd),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
defparam \Selector31~0 .lut_mask = 16'hEEFF;
defparam \Selector31~0 .sum_lutc_input = "datac";

dffeas \m_state.010000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.010000000~q ),
	.prn(vcc));
defparam \m_state.010000000 .is_wysiwyg = "true";
defparam \m_state.010000000 .power_up = "low";

cycloneive_lcell_comb \Selector35~2 (
	.dataa(\m_state.000000010~q ),
	.datab(\m_state.100000000~q ),
	.datac(\m_next~22_combout ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector35~2_combout ),
	.cout());
defparam \Selector35~2 .lut_mask = 16'hBFFF;
defparam \Selector35~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~0 (
	.dataa(\active_rnw~q ),
	.datab(\Selector35~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector34~0_combout ),
	.cout());
defparam \Selector34~0 .lut_mask = 16'hEEEE;
defparam \Selector34~0 .sum_lutc_input = "datac";

dffeas \m_next.000001000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector34~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector34~2_combout ),
	.q(\m_next.000001000~q ),
	.prn(vcc));
defparam \m_next.000001000 .is_wysiwyg = "true";
defparam \m_next.000001000 .power_up = "low";

cycloneive_lcell_comb \Selector27~2 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.datab(\m_next.000001000~q ),
	.datac(\Selector27~0_combout ),
	.datad(\Selector27~1_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
defparam \Selector27~2 .lut_mask = 16'hFFFE;
defparam \Selector27~2 .sum_lutc_input = "datac";

dffeas \m_state.000001000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector27~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector27~6_combout ),
	.q(\m_state.000001000~q ),
	.prn(vcc));
defparam \m_state.000001000 .is_wysiwyg = "true";
defparam \m_state.000001000 .power_up = "low";

cycloneive_lcell_comb \WideOr9~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\m_state.000001000~q ),
	.datad(\m_state.000010000~q ),
	.cin(gnd),
	.combout(\WideOr9~0_combout ),
	.cout());
defparam \WideOr9~0 .lut_mask = 16'h0FFF;
defparam \WideOr9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~1 (
	.dataa(\Selector32~0_combout ),
	.datab(\pending~combout ),
	.datac(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector32~1_combout ),
	.cout());
defparam \Selector32~1 .lut_mask = 16'hEFFF;
defparam \Selector32~1 .sum_lutc_input = "datac";

dffeas \m_state.100000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector32~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.100000000~q ),
	.prn(vcc));
defparam \m_state.100000000 .is_wysiwyg = "true";
defparam \m_state.100000000 .power_up = "low";

cycloneive_lcell_comb \Selector26~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_state.100000000~q ),
	.datac(\refresh_request~q ),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
defparam \Selector26~0 .lut_mask = 16'hFFFE;
defparam \Selector26~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~1 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
defparam \Selector26~1 .lut_mask = 16'hFFFE;
defparam \Selector26~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~2 (
	.dataa(\Selector26~0_combout ),
	.datab(\Selector26~1_combout ),
	.datac(\pending~combout ),
	.datad(\WideOr8~0_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
defparam \Selector26~2 .lut_mask = 16'hEFFF;
defparam \Selector26~2 .sum_lutc_input = "datac";

dffeas \m_state.000000100 (
	.clk(wire_pll7_clk_0),
	.d(\Selector26~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000100~q ),
	.prn(vcc));
defparam \m_state.000000100 .is_wysiwyg = "true";
defparam \m_state.000000100 .power_up = "low";

cycloneive_lcell_comb \Selector24~0 (
	.dataa(\m_state.000000100~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
defparam \Selector24~0 .lut_mask = 16'hAAFF;
defparam \Selector24~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~6 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\refresh_request~q ),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\Selector35~6_combout ),
	.cout());
defparam \Selector35~6 .lut_mask = 16'hFEFF;
defparam \Selector35~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector33~1_combout ),
	.cout());
defparam \Selector33~1 .lut_mask = 16'h0FFF;
defparam \Selector33~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~2 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000000001~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector33~2_combout ),
	.cout());
defparam \Selector33~2 .lut_mask = 16'hEFFF;
defparam \Selector33~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~3 (
	.dataa(\m_state.100000000~q ),
	.datab(\Selector33~2_combout ),
	.datac(\Selector33~0_combout ),
	.datad(\m_next.000000001~q ),
	.cin(gnd),
	.combout(\Selector33~3_combout ),
	.cout());
defparam \Selector33~3 .lut_mask = 16'hEFFF;
defparam \Selector33~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~4 (
	.dataa(\Selector35~6_combout ),
	.datab(\Selector33~1_combout ),
	.datac(\Selector33~3_combout ),
	.datad(\Selector35~4_combout ),
	.cin(gnd),
	.combout(\Selector33~4_combout ),
	.cout());
defparam \Selector33~4 .lut_mask = 16'hFF7F;
defparam \Selector33~4 .sum_lutc_input = "datac";

dffeas \m_next.000000001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector33~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.000000001~q ),
	.prn(vcc));
defparam \m_next.000000001 .is_wysiwyg = "true";
defparam \m_next.000000001 .power_up = "low";

cycloneive_lcell_comb \Selector24~2 (
	.dataa(\Selector24~1_combout ),
	.datab(\Selector24~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\m_next.000000001~q ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
defparam \Selector24~2 .lut_mask = 16'hFFF7;
defparam \Selector24~2 .sum_lutc_input = "datac";

dffeas \m_state.000000001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector24~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000001~q ),
	.prn(vcc));
defparam \m_state.000000001 .is_wysiwyg = "true";
defparam \m_state.000000001 .power_up = "low";

cycloneive_lcell_comb \Selector23~0 (
	.dataa(\m_state.000000001~q ),
	.datab(\ack_refresh_request~q ),
	.datac(\m_state.010000000~q ),
	.datad(\init_done~q ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
defparam \Selector23~0 .lut_mask = 16'hFEFF;
defparam \Selector23~0 .sum_lutc_input = "datac";

dffeas ack_refresh_request(
	.clk(wire_pll7_clk_0),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ack_refresh_request~q ),
	.prn(vcc));
defparam ack_refresh_request.is_wysiwyg = "true";
defparam ack_refresh_request.power_up = "low";

cycloneive_lcell_comb \refresh_request~0 (
	.dataa(\init_done~q ),
	.datab(\refresh_request~q ),
	.datac(\Equal0~4_combout ),
	.datad(\ack_refresh_request~q ),
	.cin(gnd),
	.combout(\refresh_request~0_combout ),
	.cout());
defparam \refresh_request~0 .lut_mask = 16'hFEFF;
defparam \refresh_request~0 .sum_lutc_input = "datac";

dffeas refresh_request(
	.clk(wire_pll7_clk_0),
	.d(\refresh_request~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_request~q ),
	.prn(vcc));
defparam refresh_request.is_wysiwyg = "true";
defparam refresh_request.power_up = "low";

cycloneive_lcell_comb \active_cs_n~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\init_done~q ),
	.datac(gnd),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\active_cs_n~0_combout ),
	.cout());
defparam \active_cs_n~0 .lut_mask = 16'hEEFF;
defparam \active_cs_n~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_cs_n~1 (
	.dataa(\refresh_request~q ),
	.datab(\active_cs_n~q ),
	.datac(\active_cs_n~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.cin(gnd),
	.combout(\active_cs_n~1_combout ),
	.cout());
defparam \active_cs_n~1 .lut_mask = 16'hACFF;
defparam \active_cs_n~1 .sum_lutc_input = "datac";

dffeas active_cs_n(
	.clk(wire_pll7_clk_0),
	.d(\active_cs_n~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\active_cs_n~q ),
	.prn(vcc));
defparam active_cs_n.is_wysiwyg = "true";
defparam active_cs_n.power_up = "low";

cycloneive_lcell_comb pending(
	.dataa(\active_cs_n~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\pending~4_combout ),
	.datad(\pending~9_combout ),
	.cin(gnd),
	.combout(\pending~combout ),
	.cout());
defparam pending.lut_mask = 16'hBFFF;
defparam pending.sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~2 (
	.dataa(\pending~combout ),
	.datab(\refresh_request~q ),
	.datac(\m_state.000001000~q ),
	.datad(\m_state.000010000~q ),
	.cin(gnd),
	.combout(\active_rnw~2_combout ),
	.cout());
defparam \active_rnw~2 .lut_mask = 16'hEFFF;
defparam \active_rnw~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~4 (
	.dataa(\init_done~q ),
	.datab(\m_state.000000001~q ),
	.datac(\m_state.100000000~q ),
	.datad(\Selector25~5_combout ),
	.cin(gnd),
	.combout(\active_rnw~4_combout ),
	.cout());
defparam \active_rnw~4 .lut_mask = 16'hDFFF;
defparam \active_rnw~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~3 (
	.dataa(\active_rnw~2_combout ),
	.datab(\Selector29~0_combout ),
	.datac(\active_rnw~4_combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\active_rnw~3_combout ),
	.cout());
defparam \active_rnw~3 .lut_mask = 16'hFF7F;
defparam \active_rnw~3 .sum_lutc_input = "datac";

dffeas \active_addr[11] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[47]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[11]~q ),
	.prn(vcc));
defparam \active_addr[11] .is_wysiwyg = "true";
defparam \active_addr[11] .power_up = "low";

cycloneive_lcell_comb \Selector41~0 (
	.dataa(\m_state.100000000~q ),
	.datab(entries_1),
	.datac(entries_0),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
defparam \Selector41~0 .lut_mask = 16'hFEFF;
defparam \Selector41~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector41~1 (
	.dataa(\Selector25~6_combout ),
	.datab(\pending~10_combout ),
	.datac(\Selector41~0_combout ),
	.datad(\active_rnw~2_combout ),
	.cin(gnd),
	.combout(\Selector41~1_combout ),
	.cout());
defparam \Selector41~1 .lut_mask = 16'hFEFF;
defparam \Selector41~1 .sum_lutc_input = "datac";

dffeas f_pop(
	.clk(wire_pll7_clk_0),
	.d(\Selector41~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\f_pop~q ),
	.prn(vcc));
defparam f_pop.is_wysiwyg = "true";
defparam f_pop.power_up = "low";

cycloneive_lcell_comb \m_addr[3]~0 (
	.dataa(\m_state.000000010~q ),
	.datab(\WideOr9~0_combout ),
	.datac(\f_pop~q ),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\m_addr[3]~0_combout ),
	.cout());
defparam \m_addr[3]~0 .lut_mask = 16'hB8FF;
defparam \m_addr[3]~0 .sum_lutc_input = "datac";

dffeas \active_addr[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[36]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[0]~q ),
	.prn(vcc));
defparam \active_addr[0] .is_wysiwyg = "true";
defparam \active_addr[0] .power_up = "low";

dffeas \i_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\i_state.111~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_addr[12]~q ),
	.prn(vcc));
defparam \i_addr[12] .is_wysiwyg = "true";
defparam \i_addr[12] .power_up = "low";

cycloneive_lcell_comb \Selector116~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[0]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector116~0_combout ),
	.cout());
defparam \Selector116~0 .lut_mask = 16'hDEFF;
defparam \Selector116~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector116~1 (
	.dataa(\active_addr[11]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector116~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[36]~16_combout ),
	.cin(gnd),
	.combout(\Selector116~1_combout ),
	.cout());
defparam \Selector116~1 .lut_mask = 16'hFFBE;
defparam \Selector116~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_addr[3]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\m_addr[3]~1_combout ),
	.cout());
defparam \m_addr[3]~1 .lut_mask = 16'h0FFF;
defparam \m_addr[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_addr[3]~2 (
	.dataa(\m_state.010000000~q ),
	.datab(\m_state.100000000~q ),
	.datac(\Selector25~4_combout ),
	.datad(\m_addr[3]~1_combout ),
	.cin(gnd),
	.combout(\m_addr[3]~2_combout ),
	.cout());
defparam \m_addr[3]~2 .lut_mask = 16'hFF7F;
defparam \m_addr[3]~2 .sum_lutc_input = "datac";

dffeas \active_addr[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[37]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[1]~q ),
	.prn(vcc));
defparam \active_addr[1] .is_wysiwyg = "true";
defparam \active_addr[1] .power_up = "low";

cycloneive_lcell_comb \Selector115~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[1]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector115~0_combout ),
	.cout());
defparam \Selector115~0 .lut_mask = 16'hDEFF;
defparam \Selector115~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector115~1 (
	.dataa(\active_addr[12]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector115~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[37]~17_combout ),
	.cin(gnd),
	.combout(\Selector115~1_combout ),
	.cout());
defparam \Selector115~1 .lut_mask = 16'hFFBE;
defparam \Selector115~1 .sum_lutc_input = "datac";

dffeas \active_addr[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[38]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[2]~q ),
	.prn(vcc));
defparam \active_addr[2] .is_wysiwyg = "true";
defparam \active_addr[2] .power_up = "low";

cycloneive_lcell_comb \Selector114~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[2]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector114~0_combout ),
	.cout());
defparam \Selector114~0 .lut_mask = 16'hDEFF;
defparam \Selector114~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector114~1 (
	.dataa(\active_addr[13]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector114~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[38]~18_combout ),
	.cin(gnd),
	.combout(\Selector114~1_combout ),
	.cout());
defparam \Selector114~1 .lut_mask = 16'hFFBE;
defparam \Selector114~1 .sum_lutc_input = "datac";

dffeas \active_addr[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[39]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[3]~q ),
	.prn(vcc));
defparam \active_addr[3] .is_wysiwyg = "true";
defparam \active_addr[3] .power_up = "low";

cycloneive_lcell_comb \Selector113~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[3]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector113~0_combout ),
	.cout());
defparam \Selector113~0 .lut_mask = 16'hDEFF;
defparam \Selector113~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector113~1 (
	.dataa(\active_addr[14]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector113~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[39]~19_combout ),
	.cin(gnd),
	.combout(\Selector113~1_combout ),
	.cout());
defparam \Selector113~1 .lut_mask = 16'hFFBE;
defparam \Selector113~1 .sum_lutc_input = "datac";

dffeas \active_addr[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[40]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[4]~q ),
	.prn(vcc));
defparam \active_addr[4] .is_wysiwyg = "true";
defparam \active_addr[4] .power_up = "low";

cycloneive_lcell_comb f_select(
	.dataa(\f_pop~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\f_select~combout ),
	.cout());
defparam f_select.lut_mask = 16'hAAFF;
defparam f_select.sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector112~0 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[40]~20_combout ),
	.datab(\active_addr[4]~q ),
	.datac(\f_select~combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector112~0_combout ),
	.cout());
defparam \Selector112~0 .lut_mask = 16'hACFF;
defparam \Selector112~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector112~1 (
	.dataa(\Selector112~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\active_addr[15]~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector112~1_combout ),
	.cout());
defparam \Selector112~1 .lut_mask = 16'hFEFF;
defparam \Selector112~1 .sum_lutc_input = "datac";

dffeas \active_addr[5] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[41]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[5]~q ),
	.prn(vcc));
defparam \active_addr[5] .is_wysiwyg = "true";
defparam \active_addr[5] .power_up = "low";

cycloneive_lcell_comb \Selector111~0 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[41]~21_combout ),
	.datab(\active_addr[5]~q ),
	.datac(\f_select~combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector111~0_combout ),
	.cout());
defparam \Selector111~0 .lut_mask = 16'hACFF;
defparam \Selector111~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector111~1 (
	.dataa(\Selector111~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\active_addr[16]~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector111~1_combout ),
	.cout());
defparam \Selector111~1 .lut_mask = 16'hFEFF;
defparam \Selector111~1 .sum_lutc_input = "datac";

dffeas \active_addr[6] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[42]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[6]~q ),
	.prn(vcc));
defparam \active_addr[6] .is_wysiwyg = "true";
defparam \active_addr[6] .power_up = "low";

cycloneive_lcell_comb \Selector110~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[6]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector110~0_combout ),
	.cout());
defparam \Selector110~0 .lut_mask = 16'hDEFF;
defparam \Selector110~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector110~1 (
	.dataa(\active_addr[17]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector110~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[42]~22_combout ),
	.cin(gnd),
	.combout(\Selector110~1_combout ),
	.cout());
defparam \Selector110~1 .lut_mask = 16'hFFBE;
defparam \Selector110~1 .sum_lutc_input = "datac";

dffeas \active_addr[7] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[43]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[7]~q ),
	.prn(vcc));
defparam \active_addr[7] .is_wysiwyg = "true";
defparam \active_addr[7] .power_up = "low";

cycloneive_lcell_comb \Selector109~0 (
	.dataa(\WideOr9~0_combout ),
	.datab(\active_addr[18]~q ),
	.datac(\m_addr[3]~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector109~0_combout ),
	.cout());
defparam \Selector109~0 .lut_mask = 16'hDEFF;
defparam \Selector109~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector109~1 (
	.dataa(\active_addr[7]~q ),
	.datab(\WideOr9~0_combout ),
	.datac(\Selector109~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[43]~23_combout ),
	.cin(gnd),
	.combout(\Selector109~1_combout ),
	.cout());
defparam \Selector109~1 .lut_mask = 16'hFFBE;
defparam \Selector109~1 .sum_lutc_input = "datac";

dffeas \active_addr[8] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[44]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[8]~q ),
	.prn(vcc));
defparam \active_addr[8] .is_wysiwyg = "true";
defparam \active_addr[8] .power_up = "low";

cycloneive_lcell_comb \Selector108~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[8]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector108~0_combout ),
	.cout());
defparam \Selector108~0 .lut_mask = 16'hDEFF;
defparam \Selector108~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector108~1 (
	.dataa(\active_addr[19]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector108~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[44]~24_combout ),
	.cin(gnd),
	.combout(\Selector108~1_combout ),
	.cout());
defparam \Selector108~1 .lut_mask = 16'hFFBE;
defparam \Selector108~1 .sum_lutc_input = "datac";

dffeas \active_addr[9] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[45]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[9]~q ),
	.prn(vcc));
defparam \active_addr[9] .is_wysiwyg = "true";
defparam \active_addr[9] .power_up = "low";

cycloneive_lcell_comb \Selector107~0 (
	.dataa(\WideOr9~0_combout ),
	.datab(\active_addr[20]~q ),
	.datac(\m_addr[3]~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector107~0_combout ),
	.cout());
defparam \Selector107~0 .lut_mask = 16'hDEFF;
defparam \Selector107~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector107~1 (
	.dataa(\active_addr[9]~q ),
	.datab(\WideOr9~0_combout ),
	.datac(\Selector107~0_combout ),
	.datad(\the_usb_system_sdram_input_efifo_module|rd_data[45]~25_combout ),
	.cin(gnd),
	.combout(\Selector107~1_combout ),
	.cout());
defparam \Selector107~1 .lut_mask = 16'hFFBE;
defparam \Selector107~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\pending~combout ),
	.datab(\f_pop~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'h7777;
defparam \always5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector106~2 (
	.dataa(\active_addr[21]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector106~2_combout ),
	.cout());
defparam \Selector106~2 .lut_mask = 16'h88BB;
defparam \Selector106~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector106~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector106~2_combout ),
	.cin(gnd),
	.combout(\Selector106~3_combout ),
	.cout());
defparam \Selector106~3 .lut_mask = 16'hFFF7;
defparam \Selector106~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector105~2 (
	.dataa(\active_addr[22]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector105~2_combout ),
	.cout());
defparam \Selector105~2 .lut_mask = 16'h88BB;
defparam \Selector105~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector105~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector105~2_combout ),
	.cin(gnd),
	.combout(\Selector105~3_combout ),
	.cout());
defparam \Selector105~3 .lut_mask = 16'hFFF7;
defparam \Selector105~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector104~2 (
	.dataa(\active_addr[23]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector104~2_combout ),
	.cout());
defparam \Selector104~2 .lut_mask = 16'h88BB;
defparam \Selector104~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector104~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector104~2_combout ),
	.cin(gnd),
	.combout(\Selector104~3_combout ),
	.cout());
defparam \Selector104~3 .lut_mask = 16'hFFF7;
defparam \Selector104~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector118~0 (
	.dataa(\active_addr[10]~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector118~0_combout ),
	.cout());
defparam \Selector118~0 .lut_mask = 16'hEFFE;
defparam \Selector118~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr16~0 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000000010~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr16~0_combout ),
	.cout());
defparam \WideOr16~0 .lut_mask = 16'hFEFE;
defparam \WideOr16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector117~0 (
	.dataa(\active_addr[24]~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector117~0_combout ),
	.cout());
defparam \Selector117~0 .lut_mask = 16'hEFFE;
defparam \Selector117~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\i_state.001~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[1]~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFFF7;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \i_cmd[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[1]~q ),
	.prn(vcc));
defparam \i_cmd[1] .is_wysiwyg = "true";
defparam \i_cmd[1] .power_up = "low";

cycloneive_lcell_comb \Selector21~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[1]~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
defparam \Selector21~0 .lut_mask = 16'hDFD5;
defparam \Selector21~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector21~1 (
	.dataa(\always5~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\Selector21~0_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
defparam \Selector21~1 .lut_mask = 16'hFFB8;
defparam \Selector21~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\i_state.101~q ),
	.datab(gnd),
	.datac(\i_cmd[3]~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFFF5;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \i_cmd[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[3]~q ),
	.prn(vcc));
defparam \i_cmd[3] .is_wysiwyg = "true";
defparam \i_cmd[3] .power_up = "low";

cycloneive_lcell_comb \Selector19~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[3]~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
defparam \Selector19~0 .lut_mask = 16'h27FF;
defparam \Selector19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~1 (
	.dataa(\m_state.000000001~q ),
	.datab(\m_state.001000000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
defparam \Selector19~1 .lut_mask = 16'hBFFF;
defparam \Selector19~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~2 (
	.dataa(\m_state.001000000~q ),
	.datab(\m_state.000000100~q ),
	.datac(\refresh_request~q ),
	.datad(\m_next.010000000~q ),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
defparam \Selector19~2 .lut_mask = 16'hEFFF;
defparam \Selector19~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~3 (
	.dataa(\Selector19~0_combout ),
	.datab(\active_cs_n~q ),
	.datac(\Selector19~1_combout ),
	.datad(\Selector19~2_combout ),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
defparam \Selector19~3 .lut_mask = 16'h7FFF;
defparam \Selector19~3 .sum_lutc_input = "datac";

dffeas \active_dqm[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[32]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[0]~q ),
	.prn(vcc));
defparam \active_dqm[0] .is_wysiwyg = "true";
defparam \active_dqm[0] .power_up = "low";

cycloneive_lcell_comb \Selector154~0 (
	.dataa(\active_dqm[0]~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|rd_data[32]~26_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector154~0_combout ),
	.cout());
defparam \Selector154~0 .lut_mask = 16'hEFFE;
defparam \Selector154~0 .sum_lutc_input = "datac";

dffeas \active_dqm[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[33]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[1]~q ),
	.prn(vcc));
defparam \active_dqm[1] .is_wysiwyg = "true";
defparam \active_dqm[1] .power_up = "low";

cycloneive_lcell_comb \Selector153~0 (
	.dataa(\active_dqm[1]~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|rd_data[33]~27_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector153~0_combout ),
	.cout());
defparam \Selector153~0 .lut_mask = 16'hEFFE;
defparam \Selector153~0 .sum_lutc_input = "datac";

dffeas \active_dqm[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[34]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[2]~q ),
	.prn(vcc));
defparam \active_dqm[2] .is_wysiwyg = "true";
defparam \active_dqm[2] .power_up = "low";

cycloneive_lcell_comb \Selector152~0 (
	.dataa(\active_dqm[2]~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|rd_data[34]~28_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector152~0_combout ),
	.cout());
defparam \Selector152~0 .lut_mask = 16'hEFFE;
defparam \Selector152~0 .sum_lutc_input = "datac";

dffeas \active_dqm[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[35]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[3]~q ),
	.prn(vcc));
defparam \active_dqm[3] .is_wysiwyg = "true";
defparam \active_dqm[3] .power_up = "low";

cycloneive_lcell_comb \Selector151~0 (
	.dataa(\active_dqm[3]~q ),
	.datab(\the_usb_system_sdram_input_efifo_module|rd_data[35]~29_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector151~0_combout ),
	.cout());
defparam \Selector151~0 .lut_mask = 16'hEFFE;
defparam \Selector151~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[2]~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFFF7;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \i_cmd[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[2]~q ),
	.prn(vcc));
defparam \i_cmd[2] .is_wysiwyg = "true";
defparam \i_cmd[2] .power_up = "low";

cycloneive_lcell_comb \Selector20~0 (
	.dataa(\WideOr8~0_combout ),
	.datab(\init_done~q ),
	.datac(\i_cmd[2]~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
defparam \Selector20~0 .lut_mask = 16'hF377;
defparam \Selector20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\i_state.010~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[0]~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFFF7;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \i_cmd[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[0]~q ),
	.prn(vcc));
defparam \i_cmd[0] .is_wysiwyg = "true";
defparam \i_cmd[0] .power_up = "low";

cycloneive_lcell_comb \Selector22~0 (
	.dataa(\init_done~q ),
	.datab(gnd),
	.datac(\i_cmd[0]~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
defparam \Selector22~0 .lut_mask = 16'hAFFF;
defparam \Selector22~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector22~1 (
	.dataa(\Selector22~0_combout ),
	.datab(\always5~0_combout ),
	.datac(\WideOr10~0_combout ),
	.datad(\m_state.000010000~q ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
defparam \Selector22~1 .lut_mask = 16'hCF5F;
defparam \Selector22~1 .sum_lutc_input = "datac";

dffeas \active_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[0]~q ),
	.prn(vcc));
defparam \active_data[0] .is_wysiwyg = "true";
defparam \active_data[0] .power_up = "low";

cycloneive_lcell_comb \Selector150~0 (
	.dataa(\active_data[0]~q ),
	.datab(m_data_0),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector150~0_combout ),
	.cout());
defparam \Selector150~0 .lut_mask = 16'hEFFE;
defparam \Selector150~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_data[30]~0 (
	.dataa(\f_pop~q ),
	.datab(\m_state.000010000~q ),
	.datac(gnd),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\m_data[30]~0_combout ),
	.cout());
defparam \m_data[30]~0 .lut_mask = 16'hEEFF;
defparam \m_data[30]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector150~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.datab(\Selector150~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector150~1_combout ),
	.cout());
defparam \Selector150~1 .lut_mask = 16'hAACC;
defparam \Selector150~1 .sum_lutc_input = "datac";

dffeas \active_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[1]~q ),
	.prn(vcc));
defparam \active_data[1] .is_wysiwyg = "true";
defparam \active_data[1] .power_up = "low";

cycloneive_lcell_comb \Selector149~0 (
	.dataa(\active_data[1]~q ),
	.datab(m_data_1),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector149~0_combout ),
	.cout());
defparam \Selector149~0 .lut_mask = 16'hEFFE;
defparam \Selector149~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector149~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.datab(\Selector149~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector149~1_combout ),
	.cout());
defparam \Selector149~1 .lut_mask = 16'hAACC;
defparam \Selector149~1 .sum_lutc_input = "datac";

dffeas \active_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[2]~q ),
	.prn(vcc));
defparam \active_data[2] .is_wysiwyg = "true";
defparam \active_data[2] .power_up = "low";

cycloneive_lcell_comb \Selector148~0 (
	.dataa(\active_data[2]~q ),
	.datab(m_data_2),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector148~0_combout ),
	.cout());
defparam \Selector148~0 .lut_mask = 16'hEFFE;
defparam \Selector148~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector148~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.datab(\Selector148~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector148~1_combout ),
	.cout());
defparam \Selector148~1 .lut_mask = 16'hAACC;
defparam \Selector148~1 .sum_lutc_input = "datac";

dffeas \active_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[3]~q ),
	.prn(vcc));
defparam \active_data[3] .is_wysiwyg = "true";
defparam \active_data[3] .power_up = "low";

cycloneive_lcell_comb \Selector147~0 (
	.dataa(\active_data[3]~q ),
	.datab(m_data_3),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector147~0_combout ),
	.cout());
defparam \Selector147~0 .lut_mask = 16'hEFFE;
defparam \Selector147~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector147~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.datab(\Selector147~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector147~1_combout ),
	.cout());
defparam \Selector147~1 .lut_mask = 16'hAACC;
defparam \Selector147~1 .sum_lutc_input = "datac";

dffeas \active_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[4]~q ),
	.prn(vcc));
defparam \active_data[4] .is_wysiwyg = "true";
defparam \active_data[4] .power_up = "low";

cycloneive_lcell_comb \Selector146~0 (
	.dataa(\active_data[4]~q ),
	.datab(m_data_4),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector146~0_combout ),
	.cout());
defparam \Selector146~0 .lut_mask = 16'hEFFE;
defparam \Selector146~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector146~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.datab(\Selector146~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector146~1_combout ),
	.cout());
defparam \Selector146~1 .lut_mask = 16'hAACC;
defparam \Selector146~1 .sum_lutc_input = "datac";

dffeas \active_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[5]~q ),
	.prn(vcc));
defparam \active_data[5] .is_wysiwyg = "true";
defparam \active_data[5] .power_up = "low";

cycloneive_lcell_comb \Selector145~0 (
	.dataa(\active_data[5]~q ),
	.datab(m_data_5),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector145~0_combout ),
	.cout());
defparam \Selector145~0 .lut_mask = 16'hEFFE;
defparam \Selector145~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector145~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.datab(\Selector145~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector145~1_combout ),
	.cout());
defparam \Selector145~1 .lut_mask = 16'hAACC;
defparam \Selector145~1 .sum_lutc_input = "datac";

dffeas \active_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[6]~q ),
	.prn(vcc));
defparam \active_data[6] .is_wysiwyg = "true";
defparam \active_data[6] .power_up = "low";

cycloneive_lcell_comb \Selector144~0 (
	.dataa(\active_data[6]~q ),
	.datab(m_data_6),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector144~0_combout ),
	.cout());
defparam \Selector144~0 .lut_mask = 16'hEFFE;
defparam \Selector144~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector144~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.datab(\Selector144~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector144~1_combout ),
	.cout());
defparam \Selector144~1 .lut_mask = 16'hAACC;
defparam \Selector144~1 .sum_lutc_input = "datac";

dffeas \active_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[7]~q ),
	.prn(vcc));
defparam \active_data[7] .is_wysiwyg = "true";
defparam \active_data[7] .power_up = "low";

cycloneive_lcell_comb \Selector143~0 (
	.dataa(\active_data[7]~q ),
	.datab(m_data_7),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector143~0_combout ),
	.cout());
defparam \Selector143~0 .lut_mask = 16'hEFFE;
defparam \Selector143~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector143~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.datab(\Selector143~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector143~1_combout ),
	.cout());
defparam \Selector143~1 .lut_mask = 16'hAACC;
defparam \Selector143~1 .sum_lutc_input = "datac";

dffeas \active_data[8] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[8]~q ),
	.prn(vcc));
defparam \active_data[8] .is_wysiwyg = "true";
defparam \active_data[8] .power_up = "low";

cycloneive_lcell_comb \Selector142~0 (
	.dataa(\active_data[8]~q ),
	.datab(m_data_8),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector142~0_combout ),
	.cout());
defparam \Selector142~0 .lut_mask = 16'hEFFE;
defparam \Selector142~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector142~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.datab(\Selector142~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector142~1_combout ),
	.cout());
defparam \Selector142~1 .lut_mask = 16'hAACC;
defparam \Selector142~1 .sum_lutc_input = "datac";

dffeas \active_data[9] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[9]~q ),
	.prn(vcc));
defparam \active_data[9] .is_wysiwyg = "true";
defparam \active_data[9] .power_up = "low";

cycloneive_lcell_comb \Selector141~0 (
	.dataa(\active_data[9]~q ),
	.datab(m_data_9),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector141~0_combout ),
	.cout());
defparam \Selector141~0 .lut_mask = 16'hEFFE;
defparam \Selector141~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector141~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.datab(\Selector141~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector141~1_combout ),
	.cout());
defparam \Selector141~1 .lut_mask = 16'hAACC;
defparam \Selector141~1 .sum_lutc_input = "datac";

dffeas \active_data[10] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[10]~q ),
	.prn(vcc));
defparam \active_data[10] .is_wysiwyg = "true";
defparam \active_data[10] .power_up = "low";

cycloneive_lcell_comb \Selector140~0 (
	.dataa(\active_data[10]~q ),
	.datab(m_data_10),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector140~0_combout ),
	.cout());
defparam \Selector140~0 .lut_mask = 16'hEFFE;
defparam \Selector140~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector140~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.datab(\Selector140~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector140~1_combout ),
	.cout());
defparam \Selector140~1 .lut_mask = 16'hAACC;
defparam \Selector140~1 .sum_lutc_input = "datac";

dffeas \active_data[11] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[11]~q ),
	.prn(vcc));
defparam \active_data[11] .is_wysiwyg = "true";
defparam \active_data[11] .power_up = "low";

cycloneive_lcell_comb \Selector139~0 (
	.dataa(\active_data[11]~q ),
	.datab(m_data_11),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector139~0_combout ),
	.cout());
defparam \Selector139~0 .lut_mask = 16'hEFFE;
defparam \Selector139~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector139~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.datab(\Selector139~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector139~1_combout ),
	.cout());
defparam \Selector139~1 .lut_mask = 16'hAACC;
defparam \Selector139~1 .sum_lutc_input = "datac";

dffeas \active_data[12] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[12]~q ),
	.prn(vcc));
defparam \active_data[12] .is_wysiwyg = "true";
defparam \active_data[12] .power_up = "low";

cycloneive_lcell_comb \Selector138~0 (
	.dataa(\active_data[12]~q ),
	.datab(m_data_12),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector138~0_combout ),
	.cout());
defparam \Selector138~0 .lut_mask = 16'hEFFE;
defparam \Selector138~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector138~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.datab(\Selector138~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector138~1_combout ),
	.cout());
defparam \Selector138~1 .lut_mask = 16'hAACC;
defparam \Selector138~1 .sum_lutc_input = "datac";

dffeas \active_data[13] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[13]~q ),
	.prn(vcc));
defparam \active_data[13] .is_wysiwyg = "true";
defparam \active_data[13] .power_up = "low";

cycloneive_lcell_comb \Selector137~0 (
	.dataa(\active_data[13]~q ),
	.datab(m_data_13),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector137~0_combout ),
	.cout());
defparam \Selector137~0 .lut_mask = 16'hEFFE;
defparam \Selector137~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector137~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.datab(\Selector137~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector137~1_combout ),
	.cout());
defparam \Selector137~1 .lut_mask = 16'hAACC;
defparam \Selector137~1 .sum_lutc_input = "datac";

dffeas \active_data[14] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[14]~q ),
	.prn(vcc));
defparam \active_data[14] .is_wysiwyg = "true";
defparam \active_data[14] .power_up = "low";

cycloneive_lcell_comb \Selector136~0 (
	.dataa(\active_data[14]~q ),
	.datab(m_data_14),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector136~0_combout ),
	.cout());
defparam \Selector136~0 .lut_mask = 16'hEFFE;
defparam \Selector136~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector136~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.datab(\Selector136~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector136~1_combout ),
	.cout());
defparam \Selector136~1 .lut_mask = 16'hAACC;
defparam \Selector136~1 .sum_lutc_input = "datac";

dffeas \active_data[15] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[15]~q ),
	.prn(vcc));
defparam \active_data[15] .is_wysiwyg = "true";
defparam \active_data[15] .power_up = "low";

cycloneive_lcell_comb \Selector135~0 (
	.dataa(\active_data[15]~q ),
	.datab(m_data_15),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector135~0_combout ),
	.cout());
defparam \Selector135~0 .lut_mask = 16'hEFFE;
defparam \Selector135~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector135~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.datab(\Selector135~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector135~1_combout ),
	.cout());
defparam \Selector135~1 .lut_mask = 16'hAACC;
defparam \Selector135~1 .sum_lutc_input = "datac";

dffeas \active_data[16] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[16]~q ),
	.prn(vcc));
defparam \active_data[16] .is_wysiwyg = "true";
defparam \active_data[16] .power_up = "low";

cycloneive_lcell_comb \Selector134~0 (
	.dataa(\active_data[16]~q ),
	.datab(m_data_16),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector134~0_combout ),
	.cout());
defparam \Selector134~0 .lut_mask = 16'hEFFE;
defparam \Selector134~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector134~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.datab(\Selector134~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector134~1_combout ),
	.cout());
defparam \Selector134~1 .lut_mask = 16'hAACC;
defparam \Selector134~1 .sum_lutc_input = "datac";

dffeas \active_data[17] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[17]~q ),
	.prn(vcc));
defparam \active_data[17] .is_wysiwyg = "true";
defparam \active_data[17] .power_up = "low";

cycloneive_lcell_comb \Selector133~0 (
	.dataa(\active_data[17]~q ),
	.datab(m_data_17),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector133~0_combout ),
	.cout());
defparam \Selector133~0 .lut_mask = 16'hEFFE;
defparam \Selector133~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector133~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.datab(\Selector133~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector133~1_combout ),
	.cout());
defparam \Selector133~1 .lut_mask = 16'hAACC;
defparam \Selector133~1 .sum_lutc_input = "datac";

dffeas \active_data[18] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[18]~q ),
	.prn(vcc));
defparam \active_data[18] .is_wysiwyg = "true";
defparam \active_data[18] .power_up = "low";

cycloneive_lcell_comb \Selector132~0 (
	.dataa(\active_data[18]~q ),
	.datab(m_data_18),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector132~0_combout ),
	.cout());
defparam \Selector132~0 .lut_mask = 16'hEFFE;
defparam \Selector132~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector132~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.datab(\Selector132~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector132~1_combout ),
	.cout());
defparam \Selector132~1 .lut_mask = 16'hAACC;
defparam \Selector132~1 .sum_lutc_input = "datac";

dffeas \active_data[19] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[19]~q ),
	.prn(vcc));
defparam \active_data[19] .is_wysiwyg = "true";
defparam \active_data[19] .power_up = "low";

cycloneive_lcell_comb \Selector131~0 (
	.dataa(\active_data[19]~q ),
	.datab(m_data_19),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector131~0_combout ),
	.cout());
defparam \Selector131~0 .lut_mask = 16'hEFFE;
defparam \Selector131~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector131~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.datab(\Selector131~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector131~1_combout ),
	.cout());
defparam \Selector131~1 .lut_mask = 16'hAACC;
defparam \Selector131~1 .sum_lutc_input = "datac";

dffeas \active_data[20] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[20]~q ),
	.prn(vcc));
defparam \active_data[20] .is_wysiwyg = "true";
defparam \active_data[20] .power_up = "low";

cycloneive_lcell_comb \Selector130~0 (
	.dataa(\active_data[20]~q ),
	.datab(m_data_20),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector130~0_combout ),
	.cout());
defparam \Selector130~0 .lut_mask = 16'hEFFE;
defparam \Selector130~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector130~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.datab(\Selector130~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector130~1_combout ),
	.cout());
defparam \Selector130~1 .lut_mask = 16'hAACC;
defparam \Selector130~1 .sum_lutc_input = "datac";

dffeas \active_data[21] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[21]~q ),
	.prn(vcc));
defparam \active_data[21] .is_wysiwyg = "true";
defparam \active_data[21] .power_up = "low";

cycloneive_lcell_comb \Selector129~0 (
	.dataa(\active_data[21]~q ),
	.datab(m_data_21),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector129~0_combout ),
	.cout());
defparam \Selector129~0 .lut_mask = 16'hEFFE;
defparam \Selector129~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector129~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.datab(\Selector129~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector129~1_combout ),
	.cout());
defparam \Selector129~1 .lut_mask = 16'hAACC;
defparam \Selector129~1 .sum_lutc_input = "datac";

dffeas \active_data[22] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[22]~q ),
	.prn(vcc));
defparam \active_data[22] .is_wysiwyg = "true";
defparam \active_data[22] .power_up = "low";

cycloneive_lcell_comb \Selector128~0 (
	.dataa(\active_data[22]~q ),
	.datab(m_data_22),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector128~0_combout ),
	.cout());
defparam \Selector128~0 .lut_mask = 16'hEFFE;
defparam \Selector128~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector128~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.datab(\Selector128~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector128~1_combout ),
	.cout());
defparam \Selector128~1 .lut_mask = 16'hAACC;
defparam \Selector128~1 .sum_lutc_input = "datac";

dffeas \active_data[23] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[23]~q ),
	.prn(vcc));
defparam \active_data[23] .is_wysiwyg = "true";
defparam \active_data[23] .power_up = "low";

cycloneive_lcell_comb \Selector127~0 (
	.dataa(\active_data[23]~q ),
	.datab(m_data_23),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector127~0_combout ),
	.cout());
defparam \Selector127~0 .lut_mask = 16'hEFFE;
defparam \Selector127~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector127~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.datab(\Selector127~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector127~1_combout ),
	.cout());
defparam \Selector127~1 .lut_mask = 16'hAACC;
defparam \Selector127~1 .sum_lutc_input = "datac";

dffeas \active_data[24] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[24]~q ),
	.prn(vcc));
defparam \active_data[24] .is_wysiwyg = "true";
defparam \active_data[24] .power_up = "low";

cycloneive_lcell_comb \Selector126~0 (
	.dataa(\active_data[24]~q ),
	.datab(m_data_24),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector126~0_combout ),
	.cout());
defparam \Selector126~0 .lut_mask = 16'hEFFE;
defparam \Selector126~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector126~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.datab(\Selector126~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector126~1_combout ),
	.cout());
defparam \Selector126~1 .lut_mask = 16'hAACC;
defparam \Selector126~1 .sum_lutc_input = "datac";

dffeas \active_data[25] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[25]~q ),
	.prn(vcc));
defparam \active_data[25] .is_wysiwyg = "true";
defparam \active_data[25] .power_up = "low";

cycloneive_lcell_comb \Selector125~0 (
	.dataa(\active_data[25]~q ),
	.datab(m_data_25),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector125~0_combout ),
	.cout());
defparam \Selector125~0 .lut_mask = 16'hEFFE;
defparam \Selector125~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector125~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.datab(\Selector125~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector125~1_combout ),
	.cout());
defparam \Selector125~1 .lut_mask = 16'hAACC;
defparam \Selector125~1 .sum_lutc_input = "datac";

dffeas \active_data[26] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[26]~q ),
	.prn(vcc));
defparam \active_data[26] .is_wysiwyg = "true";
defparam \active_data[26] .power_up = "low";

cycloneive_lcell_comb \Selector124~0 (
	.dataa(\active_data[26]~q ),
	.datab(m_data_26),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector124~0_combout ),
	.cout());
defparam \Selector124~0 .lut_mask = 16'hEFFE;
defparam \Selector124~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector124~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.datab(\Selector124~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector124~1_combout ),
	.cout());
defparam \Selector124~1 .lut_mask = 16'hAACC;
defparam \Selector124~1 .sum_lutc_input = "datac";

dffeas \active_data[27] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[27]~q ),
	.prn(vcc));
defparam \active_data[27] .is_wysiwyg = "true";
defparam \active_data[27] .power_up = "low";

cycloneive_lcell_comb \Selector123~0 (
	.dataa(\active_data[27]~q ),
	.datab(m_data_27),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector123~0_combout ),
	.cout());
defparam \Selector123~0 .lut_mask = 16'hEFFE;
defparam \Selector123~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector123~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.datab(\Selector123~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector123~1_combout ),
	.cout());
defparam \Selector123~1 .lut_mask = 16'hAACC;
defparam \Selector123~1 .sum_lutc_input = "datac";

dffeas \active_data[28] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[28]~q ),
	.prn(vcc));
defparam \active_data[28] .is_wysiwyg = "true";
defparam \active_data[28] .power_up = "low";

cycloneive_lcell_comb \Selector122~0 (
	.dataa(\active_data[28]~q ),
	.datab(m_data_28),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector122~0_combout ),
	.cout());
defparam \Selector122~0 .lut_mask = 16'hEFFE;
defparam \Selector122~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector122~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.datab(\Selector122~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector122~1_combout ),
	.cout());
defparam \Selector122~1 .lut_mask = 16'hAACC;
defparam \Selector122~1 .sum_lutc_input = "datac";

dffeas \active_data[29] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[29]~q ),
	.prn(vcc));
defparam \active_data[29] .is_wysiwyg = "true";
defparam \active_data[29] .power_up = "low";

cycloneive_lcell_comb \Selector121~0 (
	.dataa(\active_data[29]~q ),
	.datab(m_data_29),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector121~0_combout ),
	.cout());
defparam \Selector121~0 .lut_mask = 16'hEFFE;
defparam \Selector121~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector121~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.datab(\Selector121~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector121~1_combout ),
	.cout());
defparam \Selector121~1 .lut_mask = 16'hAACC;
defparam \Selector121~1 .sum_lutc_input = "datac";

dffeas \active_data[30] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[30]~q ),
	.prn(vcc));
defparam \active_data[30] .is_wysiwyg = "true";
defparam \active_data[30] .power_up = "low";

cycloneive_lcell_comb \Selector120~0 (
	.dataa(\active_data[30]~q ),
	.datab(m_data_30),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector120~0_combout ),
	.cout());
defparam \Selector120~0 .lut_mask = 16'hEFFE;
defparam \Selector120~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector120~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.datab(\Selector120~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector120~1_combout ),
	.cout());
defparam \Selector120~1 .lut_mask = 16'hAACC;
defparam \Selector120~1 .sum_lutc_input = "datac";

dffeas \active_data[31] (
	.clk(wire_pll7_clk_0),
	.d(\the_usb_system_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[31]~q ),
	.prn(vcc));
defparam \active_data[31] .is_wysiwyg = "true";
defparam \active_data[31] .power_up = "low";

cycloneive_lcell_comb \Selector119~0 (
	.dataa(\active_data[31]~q ),
	.datab(m_data_31),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector119~0_combout ),
	.cout());
defparam \Selector119~0 .lut_mask = 16'hEFFE;
defparam \Selector119~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector119~1 (
	.dataa(\the_usb_system_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.datab(\Selector119~0_combout ),
	.datac(gnd),
	.datad(\m_data[30]~0_combout ),
	.cin(gnd),
	.combout(\Selector119~1_combout ),
	.cout());
defparam \Selector119~1 .lut_mask = 16'hAACC;
defparam \Selector119~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~0 (
	.dataa(m_cmd_1),
	.datab(gnd),
	.datac(m_cmd_2),
	.datad(m_cmd_0),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hAFFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

dffeas \rd_valid[0] (
	.clk(wire_pll7_clk_0),
	.d(\Equal4~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[0]~q ),
	.prn(vcc));
defparam \rd_valid[0] .is_wysiwyg = "true";
defparam \rd_valid[0] .power_up = "low";

dffeas \rd_valid[1] (
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[1]~q ),
	.prn(vcc));
defparam \rd_valid[1] .is_wysiwyg = "true";
defparam \rd_valid[1] .power_up = "low";

dffeas \rd_valid[2] (
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[2]~q ),
	.prn(vcc));
defparam \rd_valid[2] .is_wysiwyg = "true";
defparam \rd_valid[2] .power_up = "low";

endmodule

module usb_system_usb_system_sdram_input_efifo_module (
	clk,
	f_pop,
	entries_1,
	entries_0,
	Equal1,
	rd_data_46,
	rd_data_61,
	rd_data_60,
	rd_data_47,
	rd_data_49,
	rd_data_48,
	rd_data_51,
	rd_data_50,
	rd_data_53,
	rd_data_52,
	rd_data_55,
	rd_data_54,
	rd_data_57,
	rd_data_56,
	rd_data_59,
	rd_data_58,
	pending,
	rd_data_36,
	reset_n,
	rd_data_37,
	rd_data_38,
	rd_data_39,
	rd_data_40,
	f_select,
	rd_data_41,
	rd_data_42,
	rd_data_43,
	rd_data_44,
	rd_data_45,
	rd_data_32,
	rd_data_33,
	rd_data_34,
	rd_data_35,
	last_cycle,
	WideOr1,
	src_payload,
	src_data_68,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	src_data_61,
	src_data_60,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	comb,
	comb1,
	comb2,
	comb3,
	rd_data_0,
	rd_data_1,
	rd_data_2,
	rd_data_3,
	rd_data_4,
	rd_data_5,
	rd_data_6,
	rd_data_7,
	rd_data_8,
	rd_data_9,
	rd_data_10,
	rd_data_11,
	rd_data_12,
	rd_data_13,
	rd_data_14,
	rd_data_15,
	rd_data_16,
	rd_data_17,
	rd_data_18,
	rd_data_19,
	rd_data_20,
	rd_data_21,
	rd_data_22,
	rd_data_23,
	rd_data_24,
	rd_data_25,
	rd_data_26,
	rd_data_27,
	rd_data_28,
	rd_data_29,
	rd_data_30,
	rd_data_31,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	f_pop;
output 	entries_1;
output 	entries_0;
output 	Equal1;
output 	rd_data_46;
output 	rd_data_61;
output 	rd_data_60;
output 	rd_data_47;
output 	rd_data_49;
output 	rd_data_48;
output 	rd_data_51;
output 	rd_data_50;
output 	rd_data_53;
output 	rd_data_52;
output 	rd_data_55;
output 	rd_data_54;
output 	rd_data_57;
output 	rd_data_56;
output 	rd_data_59;
output 	rd_data_58;
input 	pending;
output 	rd_data_36;
input 	reset_n;
output 	rd_data_37;
output 	rd_data_38;
output 	rd_data_39;
output 	rd_data_40;
input 	f_select;
output 	rd_data_41;
output 	rd_data_42;
output 	rd_data_43;
output 	rd_data_44;
output 	rd_data_45;
output 	rd_data_32;
output 	rd_data_33;
output 	rd_data_34;
output 	rd_data_35;
input 	last_cycle;
input 	WideOr1;
input 	src_payload;
input 	src_data_68;
input 	src_data_48;
input 	src_data_62;
input 	src_data_49;
input 	src_data_51;
input 	src_data_50;
input 	src_data_53;
input 	src_data_52;
input 	src_data_55;
input 	src_data_54;
input 	src_data_57;
input 	src_data_56;
input 	src_data_59;
input 	src_data_58;
input 	src_data_61;
input 	src_data_60;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	comb;
input 	comb1;
input 	comb2;
input 	comb3;
output 	rd_data_0;
output 	rd_data_1;
output 	rd_data_2;
output 	rd_data_3;
output 	rd_data_4;
output 	rd_data_5;
output 	rd_data_6;
output 	rd_data_7;
output 	rd_data_8;
output 	rd_data_9;
output 	rd_data_10;
output 	rd_data_11;
output 	rd_data_12;
output 	rd_data_13;
output 	rd_data_14;
output 	rd_data_15;
output 	rd_data_16;
output 	rd_data_17;
output 	rd_data_18;
output 	rd_data_19;
output 	rd_data_20;
output 	rd_data_21;
output 	rd_data_22;
output 	rd_data_23;
output 	rd_data_24;
output 	rd_data_25;
output 	rd_data_26;
output 	rd_data_27;
output 	rd_data_28;
output 	rd_data_29;
output 	rd_data_30;
output 	rd_data_31;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always2~0_combout ;
wire \entries[1]~0_combout ;
wire \entries[0]~1_combout ;
wire \wr_address~0_combout ;
wire \wr_address~q ;
wire \entry_1[61]~0_combout ;
wire \entry_1[46]~q ;
wire \entry_0[61]~0_combout ;
wire \entry_0[46]~q ;
wire \rd_address~0_combout ;
wire \rd_address~q ;
wire \entry_1[61]~q ;
wire \entry_0[61]~q ;
wire \entry_1[60]~q ;
wire \entry_0[60]~q ;
wire \entry_1[47]~q ;
wire \entry_0[47]~q ;
wire \entry_1[49]~q ;
wire \entry_0[49]~q ;
wire \entry_1[48]~q ;
wire \entry_0[48]~q ;
wire \entry_1[51]~q ;
wire \entry_0[51]~q ;
wire \entry_1[50]~q ;
wire \entry_0[50]~q ;
wire \entry_1[53]~q ;
wire \entry_0[53]~q ;
wire \entry_1[52]~q ;
wire \entry_0[52]~q ;
wire \entry_1[55]~q ;
wire \entry_0[55]~q ;
wire \entry_1[54]~q ;
wire \entry_0[54]~q ;
wire \entry_1[57]~q ;
wire \entry_0[57]~q ;
wire \entry_1[56]~q ;
wire \entry_0[56]~q ;
wire \entry_1[59]~q ;
wire \entry_0[59]~q ;
wire \entry_1[58]~q ;
wire \entry_0[58]~q ;
wire \entry_1[36]~q ;
wire \entry_0[36]~q ;
wire \entry_1[37]~q ;
wire \entry_0[37]~q ;
wire \entry_1[38]~q ;
wire \entry_0[38]~q ;
wire \entry_1[39]~q ;
wire \entry_0[39]~q ;
wire \entry_1[40]~q ;
wire \entry_0[40]~q ;
wire \entry_1[41]~q ;
wire \entry_0[41]~q ;
wire \entry_1[42]~q ;
wire \entry_0[42]~q ;
wire \entry_1[43]~q ;
wire \entry_0[43]~q ;
wire \entry_1[44]~q ;
wire \entry_0[44]~q ;
wire \entry_1[45]~q ;
wire \entry_0[45]~q ;
wire \entry_1[32]~q ;
wire \entry_0[32]~q ;
wire \entry_1[33]~q ;
wire \entry_0[33]~q ;
wire \entry_1[34]~q ;
wire \entry_0[34]~q ;
wire \entry_1[35]~q ;
wire \entry_0[35]~q ;
wire \entry_1[0]~q ;
wire \entry_0[0]~q ;
wire \entry_1[1]~q ;
wire \entry_0[1]~q ;
wire \entry_1[2]~q ;
wire \entry_0[2]~q ;
wire \entry_1[3]~q ;
wire \entry_0[3]~q ;
wire \entry_1[4]~q ;
wire \entry_0[4]~q ;
wire \entry_1[5]~q ;
wire \entry_0[5]~q ;
wire \entry_1[6]~q ;
wire \entry_0[6]~q ;
wire \entry_1[7]~q ;
wire \entry_0[7]~q ;
wire \entry_1[8]~q ;
wire \entry_0[8]~q ;
wire \entry_1[9]~q ;
wire \entry_0[9]~q ;
wire \entry_1[10]~q ;
wire \entry_0[10]~q ;
wire \entry_1[11]~q ;
wire \entry_0[11]~q ;
wire \entry_1[12]~q ;
wire \entry_0[12]~q ;
wire \entry_1[13]~q ;
wire \entry_0[13]~q ;
wire \entry_1[14]~q ;
wire \entry_0[14]~q ;
wire \entry_1[15]~q ;
wire \entry_0[15]~q ;
wire \entry_1[16]~q ;
wire \entry_0[16]~q ;
wire \entry_1[17]~q ;
wire \entry_0[17]~q ;
wire \entry_1[18]~q ;
wire \entry_0[18]~q ;
wire \entry_1[19]~q ;
wire \entry_0[19]~q ;
wire \entry_1[20]~q ;
wire \entry_0[20]~q ;
wire \entry_1[21]~q ;
wire \entry_0[21]~q ;
wire \entry_1[22]~q ;
wire \entry_0[22]~q ;
wire \entry_1[23]~q ;
wire \entry_0[23]~q ;
wire \entry_1[24]~q ;
wire \entry_0[24]~q ;
wire \entry_1[25]~q ;
wire \entry_0[25]~q ;
wire \entry_1[26]~q ;
wire \entry_0[26]~q ;
wire \entry_1[27]~q ;
wire \entry_0[27]~q ;
wire \entry_1[28]~q ;
wire \entry_0[28]~q ;
wire \entry_1[29]~q ;
wire \entry_0[29]~q ;
wire \entry_1[30]~q ;
wire \entry_0[30]~q ;
wire \entry_1[31]~q ;
wire \entry_0[31]~q ;


dffeas \entries[1] (
	.clk(clk),
	.d(\entries[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_1),
	.prn(vcc));
defparam \entries[1] .is_wysiwyg = "true";
defparam \entries[1] .power_up = "low";

dffeas \entries[0] (
	.clk(clk),
	.d(\entries[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_0),
	.prn(vcc));
defparam \entries[0] .is_wysiwyg = "true";
defparam \entries[0] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEEEE;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[46]~0 (
	.dataa(\entry_1[46]~q ),
	.datab(\entry_0[46]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_46),
	.cout());
defparam \rd_data[46]~0 .lut_mask = 16'hAACC;
defparam \rd_data[46]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[61]~1 (
	.dataa(\entry_1[61]~q ),
	.datab(\entry_0[61]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_61),
	.cout());
defparam \rd_data[61]~1 .lut_mask = 16'hAACC;
defparam \rd_data[61]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[60]~2 (
	.dataa(\entry_1[60]~q ),
	.datab(\entry_0[60]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_60),
	.cout());
defparam \rd_data[60]~2 .lut_mask = 16'hAACC;
defparam \rd_data[60]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[47]~3 (
	.dataa(\entry_1[47]~q ),
	.datab(\entry_0[47]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_47),
	.cout());
defparam \rd_data[47]~3 .lut_mask = 16'hAACC;
defparam \rd_data[47]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[49]~4 (
	.dataa(\entry_1[49]~q ),
	.datab(\entry_0[49]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_49),
	.cout());
defparam \rd_data[49]~4 .lut_mask = 16'hAACC;
defparam \rd_data[49]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[48]~5 (
	.dataa(\entry_1[48]~q ),
	.datab(\entry_0[48]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_48),
	.cout());
defparam \rd_data[48]~5 .lut_mask = 16'hAACC;
defparam \rd_data[48]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[51]~6 (
	.dataa(\entry_1[51]~q ),
	.datab(\entry_0[51]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_51),
	.cout());
defparam \rd_data[51]~6 .lut_mask = 16'hAACC;
defparam \rd_data[51]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[50]~7 (
	.dataa(\entry_1[50]~q ),
	.datab(\entry_0[50]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_50),
	.cout());
defparam \rd_data[50]~7 .lut_mask = 16'hAACC;
defparam \rd_data[50]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[53]~8 (
	.dataa(\entry_1[53]~q ),
	.datab(\entry_0[53]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_53),
	.cout());
defparam \rd_data[53]~8 .lut_mask = 16'hAACC;
defparam \rd_data[53]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[52]~9 (
	.dataa(\entry_1[52]~q ),
	.datab(\entry_0[52]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_52),
	.cout());
defparam \rd_data[52]~9 .lut_mask = 16'hAACC;
defparam \rd_data[52]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[55]~10 (
	.dataa(\entry_1[55]~q ),
	.datab(\entry_0[55]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_55),
	.cout());
defparam \rd_data[55]~10 .lut_mask = 16'hAACC;
defparam \rd_data[55]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[54]~11 (
	.dataa(\entry_1[54]~q ),
	.datab(\entry_0[54]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_54),
	.cout());
defparam \rd_data[54]~11 .lut_mask = 16'hAACC;
defparam \rd_data[54]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[57]~12 (
	.dataa(\entry_1[57]~q ),
	.datab(\entry_0[57]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_57),
	.cout());
defparam \rd_data[57]~12 .lut_mask = 16'hAACC;
defparam \rd_data[57]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[56]~13 (
	.dataa(\entry_1[56]~q ),
	.datab(\entry_0[56]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_56),
	.cout());
defparam \rd_data[56]~13 .lut_mask = 16'hAACC;
defparam \rd_data[56]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[59]~14 (
	.dataa(\entry_1[59]~q ),
	.datab(\entry_0[59]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_59),
	.cout());
defparam \rd_data[59]~14 .lut_mask = 16'hAACC;
defparam \rd_data[59]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[58]~15 (
	.dataa(\entry_1[58]~q ),
	.datab(\entry_0[58]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_58),
	.cout());
defparam \rd_data[58]~15 .lut_mask = 16'hAACC;
defparam \rd_data[58]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[36]~16 (
	.dataa(\entry_1[36]~q ),
	.datab(\entry_0[36]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_36),
	.cout());
defparam \rd_data[36]~16 .lut_mask = 16'hAACC;
defparam \rd_data[36]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[37]~17 (
	.dataa(\entry_1[37]~q ),
	.datab(\entry_0[37]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_37),
	.cout());
defparam \rd_data[37]~17 .lut_mask = 16'hAACC;
defparam \rd_data[37]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[38]~18 (
	.dataa(\entry_1[38]~q ),
	.datab(\entry_0[38]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_38),
	.cout());
defparam \rd_data[38]~18 .lut_mask = 16'hAACC;
defparam \rd_data[38]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[39]~19 (
	.dataa(\entry_1[39]~q ),
	.datab(\entry_0[39]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_39),
	.cout());
defparam \rd_data[39]~19 .lut_mask = 16'hAACC;
defparam \rd_data[39]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[40]~20 (
	.dataa(\entry_1[40]~q ),
	.datab(\entry_0[40]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_40),
	.cout());
defparam \rd_data[40]~20 .lut_mask = 16'hAACC;
defparam \rd_data[40]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[41]~21 (
	.dataa(\entry_1[41]~q ),
	.datab(\entry_0[41]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_41),
	.cout());
defparam \rd_data[41]~21 .lut_mask = 16'hAACC;
defparam \rd_data[41]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[42]~22 (
	.dataa(\entry_1[42]~q ),
	.datab(\entry_0[42]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_42),
	.cout());
defparam \rd_data[42]~22 .lut_mask = 16'hAACC;
defparam \rd_data[42]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[43]~23 (
	.dataa(\entry_1[43]~q ),
	.datab(\entry_0[43]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_43),
	.cout());
defparam \rd_data[43]~23 .lut_mask = 16'hAACC;
defparam \rd_data[43]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[44]~24 (
	.dataa(\entry_1[44]~q ),
	.datab(\entry_0[44]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_44),
	.cout());
defparam \rd_data[44]~24 .lut_mask = 16'hAACC;
defparam \rd_data[44]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[45]~25 (
	.dataa(\entry_1[45]~q ),
	.datab(\entry_0[45]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_45),
	.cout());
defparam \rd_data[45]~25 .lut_mask = 16'hAACC;
defparam \rd_data[45]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[32]~26 (
	.dataa(\entry_1[32]~q ),
	.datab(\entry_0[32]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_32),
	.cout());
defparam \rd_data[32]~26 .lut_mask = 16'hAACC;
defparam \rd_data[32]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[33]~27 (
	.dataa(\entry_1[33]~q ),
	.datab(\entry_0[33]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_33),
	.cout());
defparam \rd_data[33]~27 .lut_mask = 16'hAACC;
defparam \rd_data[33]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[34]~28 (
	.dataa(\entry_1[34]~q ),
	.datab(\entry_0[34]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_34),
	.cout());
defparam \rd_data[34]~28 .lut_mask = 16'hAACC;
defparam \rd_data[34]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[35]~29 (
	.dataa(\entry_1[35]~q ),
	.datab(\entry_0[35]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_35),
	.cout());
defparam \rd_data[35]~29 .lut_mask = 16'hAACC;
defparam \rd_data[35]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[0]~30 (
	.dataa(\entry_1[0]~q ),
	.datab(\entry_0[0]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_0),
	.cout());
defparam \rd_data[0]~30 .lut_mask = 16'hAACC;
defparam \rd_data[0]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[1]~31 (
	.dataa(\entry_1[1]~q ),
	.datab(\entry_0[1]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_1),
	.cout());
defparam \rd_data[1]~31 .lut_mask = 16'hAACC;
defparam \rd_data[1]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[2]~32 (
	.dataa(\entry_1[2]~q ),
	.datab(\entry_0[2]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_2),
	.cout());
defparam \rd_data[2]~32 .lut_mask = 16'hAACC;
defparam \rd_data[2]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[3]~33 (
	.dataa(\entry_1[3]~q ),
	.datab(\entry_0[3]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_3),
	.cout());
defparam \rd_data[3]~33 .lut_mask = 16'hAACC;
defparam \rd_data[3]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[4]~34 (
	.dataa(\entry_1[4]~q ),
	.datab(\entry_0[4]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_4),
	.cout());
defparam \rd_data[4]~34 .lut_mask = 16'hAACC;
defparam \rd_data[4]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[5]~35 (
	.dataa(\entry_1[5]~q ),
	.datab(\entry_0[5]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_5),
	.cout());
defparam \rd_data[5]~35 .lut_mask = 16'hAACC;
defparam \rd_data[5]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[6]~36 (
	.dataa(\entry_1[6]~q ),
	.datab(\entry_0[6]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_6),
	.cout());
defparam \rd_data[6]~36 .lut_mask = 16'hAACC;
defparam \rd_data[6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[7]~37 (
	.dataa(\entry_1[7]~q ),
	.datab(\entry_0[7]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_7),
	.cout());
defparam \rd_data[7]~37 .lut_mask = 16'hAACC;
defparam \rd_data[7]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[8]~38 (
	.dataa(\entry_1[8]~q ),
	.datab(\entry_0[8]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_8),
	.cout());
defparam \rd_data[8]~38 .lut_mask = 16'hAACC;
defparam \rd_data[8]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[9]~39 (
	.dataa(\entry_1[9]~q ),
	.datab(\entry_0[9]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_9),
	.cout());
defparam \rd_data[9]~39 .lut_mask = 16'hAACC;
defparam \rd_data[9]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[10]~40 (
	.dataa(\entry_1[10]~q ),
	.datab(\entry_0[10]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_10),
	.cout());
defparam \rd_data[10]~40 .lut_mask = 16'hAACC;
defparam \rd_data[10]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[11]~41 (
	.dataa(\entry_1[11]~q ),
	.datab(\entry_0[11]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_11),
	.cout());
defparam \rd_data[11]~41 .lut_mask = 16'hAACC;
defparam \rd_data[11]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[12]~42 (
	.dataa(\entry_1[12]~q ),
	.datab(\entry_0[12]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_12),
	.cout());
defparam \rd_data[12]~42 .lut_mask = 16'hAACC;
defparam \rd_data[12]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[13]~43 (
	.dataa(\entry_1[13]~q ),
	.datab(\entry_0[13]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_13),
	.cout());
defparam \rd_data[13]~43 .lut_mask = 16'hAACC;
defparam \rd_data[13]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[14]~44 (
	.dataa(\entry_1[14]~q ),
	.datab(\entry_0[14]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_14),
	.cout());
defparam \rd_data[14]~44 .lut_mask = 16'hAACC;
defparam \rd_data[14]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[15]~45 (
	.dataa(\entry_1[15]~q ),
	.datab(\entry_0[15]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_15),
	.cout());
defparam \rd_data[15]~45 .lut_mask = 16'hAACC;
defparam \rd_data[15]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[16]~46 (
	.dataa(\entry_1[16]~q ),
	.datab(\entry_0[16]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_16),
	.cout());
defparam \rd_data[16]~46 .lut_mask = 16'hAACC;
defparam \rd_data[16]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[17]~47 (
	.dataa(\entry_1[17]~q ),
	.datab(\entry_0[17]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_17),
	.cout());
defparam \rd_data[17]~47 .lut_mask = 16'hAACC;
defparam \rd_data[17]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[18]~48 (
	.dataa(\entry_1[18]~q ),
	.datab(\entry_0[18]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_18),
	.cout());
defparam \rd_data[18]~48 .lut_mask = 16'hAACC;
defparam \rd_data[18]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[19]~49 (
	.dataa(\entry_1[19]~q ),
	.datab(\entry_0[19]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_19),
	.cout());
defparam \rd_data[19]~49 .lut_mask = 16'hAACC;
defparam \rd_data[19]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[20]~50 (
	.dataa(\entry_1[20]~q ),
	.datab(\entry_0[20]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_20),
	.cout());
defparam \rd_data[20]~50 .lut_mask = 16'hAACC;
defparam \rd_data[20]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[21]~51 (
	.dataa(\entry_1[21]~q ),
	.datab(\entry_0[21]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_21),
	.cout());
defparam \rd_data[21]~51 .lut_mask = 16'hAACC;
defparam \rd_data[21]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[22]~52 (
	.dataa(\entry_1[22]~q ),
	.datab(\entry_0[22]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_22),
	.cout());
defparam \rd_data[22]~52 .lut_mask = 16'hAACC;
defparam \rd_data[22]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[23]~53 (
	.dataa(\entry_1[23]~q ),
	.datab(\entry_0[23]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_23),
	.cout());
defparam \rd_data[23]~53 .lut_mask = 16'hAACC;
defparam \rd_data[23]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[24]~54 (
	.dataa(\entry_1[24]~q ),
	.datab(\entry_0[24]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_24),
	.cout());
defparam \rd_data[24]~54 .lut_mask = 16'hAACC;
defparam \rd_data[24]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[25]~55 (
	.dataa(\entry_1[25]~q ),
	.datab(\entry_0[25]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_25),
	.cout());
defparam \rd_data[25]~55 .lut_mask = 16'hAACC;
defparam \rd_data[25]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[26]~56 (
	.dataa(\entry_1[26]~q ),
	.datab(\entry_0[26]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_26),
	.cout());
defparam \rd_data[26]~56 .lut_mask = 16'hAACC;
defparam \rd_data[26]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[27]~57 (
	.dataa(\entry_1[27]~q ),
	.datab(\entry_0[27]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_27),
	.cout());
defparam \rd_data[27]~57 .lut_mask = 16'hAACC;
defparam \rd_data[27]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[28]~58 (
	.dataa(\entry_1[28]~q ),
	.datab(\entry_0[28]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_28),
	.cout());
defparam \rd_data[28]~58 .lut_mask = 16'hAACC;
defparam \rd_data[28]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[29]~59 (
	.dataa(\entry_1[29]~q ),
	.datab(\entry_0[29]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_29),
	.cout());
defparam \rd_data[29]~59 .lut_mask = 16'hAACC;
defparam \rd_data[29]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[30]~60 (
	.dataa(\entry_1[30]~q ),
	.datab(\entry_0[30]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_30),
	.cout());
defparam \rd_data[30]~60 .lut_mask = 16'hAACC;
defparam \rd_data[30]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[31]~61 (
	.dataa(\entry_1[31]~q ),
	.datab(\entry_0[31]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_31),
	.cout());
defparam \rd_data[31]~61 .lut_mask = 16'hAACC;
defparam \rd_data[31]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(last_cycle),
	.datab(WideOr1),
	.datac(src_payload),
	.datad(src_data_68),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hFFFE;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entries[1]~0 (
	.dataa(entries_1),
	.datab(f_select),
	.datac(entries_0),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\entries[1]~0_combout ),
	.cout());
defparam \entries[1]~0 .lut_mask = 16'h6996;
defparam \entries[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entries[0]~1 (
	.dataa(f_pop),
	.datab(pending),
	.datac(entries_0),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\entries[0]~1_combout ),
	.cout());
defparam \entries[0]~1 .lut_mask = 16'h6996;
defparam \entries[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\always2~0_combout ),
	.datad(\wr_address~q ),
	.cin(gnd),
	.combout(\wr_address~0_combout ),
	.cout());
defparam \wr_address~0 .lut_mask = 16'h0FF0;
defparam \wr_address~0 .sum_lutc_input = "datac";

dffeas wr_address(
	.clk(clk),
	.d(\wr_address~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_address~q ),
	.prn(vcc));
defparam wr_address.is_wysiwyg = "true";
defparam wr_address.power_up = "low";

cycloneive_lcell_comb \entry_1[61]~0 (
	.dataa(\always2~0_combout ),
	.datab(\wr_address~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\entry_1[61]~0_combout ),
	.cout());
defparam \entry_1[61]~0 .lut_mask = 16'hEEEE;
defparam \entry_1[61]~0 .sum_lutc_input = "datac";

dffeas \entry_1[46] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[46]~q ),
	.prn(vcc));
defparam \entry_1[46] .is_wysiwyg = "true";
defparam \entry_1[46] .power_up = "low";

cycloneive_lcell_comb \entry_0[61]~0 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wr_address~q ),
	.cin(gnd),
	.combout(\entry_0[61]~0_combout ),
	.cout());
defparam \entry_0[61]~0 .lut_mask = 16'hAAFF;
defparam \entry_0[61]~0 .sum_lutc_input = "datac";

dffeas \entry_0[46] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[46]~q ),
	.prn(vcc));
defparam \entry_0[46] .is_wysiwyg = "true";
defparam \entry_0[46] .power_up = "low";

cycloneive_lcell_comb \rd_address~0 (
	.dataa(\rd_address~q ),
	.datab(pending),
	.datac(gnd),
	.datad(f_pop),
	.cin(gnd),
	.combout(\rd_address~0_combout ),
	.cout());
defparam \rd_address~0 .lut_mask = 16'h9966;
defparam \rd_address~0 .sum_lutc_input = "datac";

dffeas rd_address(
	.clk(clk),
	.d(\rd_address~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_address~q ),
	.prn(vcc));
defparam rd_address.is_wysiwyg = "true";
defparam rd_address.power_up = "low";

dffeas \entry_1[61] (
	.clk(clk),
	.d(m0_write),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[61]~q ),
	.prn(vcc));
defparam \entry_1[61] .is_wysiwyg = "true";
defparam \entry_1[61] .power_up = "low";

dffeas \entry_0[61] (
	.clk(clk),
	.d(m0_write),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[61]~q ),
	.prn(vcc));
defparam \entry_0[61] .is_wysiwyg = "true";
defparam \entry_0[61] .power_up = "low";

dffeas \entry_1[60] (
	.clk(clk),
	.d(src_data_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[60]~q ),
	.prn(vcc));
defparam \entry_1[60] .is_wysiwyg = "true";
defparam \entry_1[60] .power_up = "low";

dffeas \entry_0[60] (
	.clk(clk),
	.d(src_data_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[60]~q ),
	.prn(vcc));
defparam \entry_0[60] .is_wysiwyg = "true";
defparam \entry_0[60] .power_up = "low";

dffeas \entry_1[47] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[47]~q ),
	.prn(vcc));
defparam \entry_1[47] .is_wysiwyg = "true";
defparam \entry_1[47] .power_up = "low";

dffeas \entry_0[47] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[47]~q ),
	.prn(vcc));
defparam \entry_0[47] .is_wysiwyg = "true";
defparam \entry_0[47] .power_up = "low";

dffeas \entry_1[49] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[49]~q ),
	.prn(vcc));
defparam \entry_1[49] .is_wysiwyg = "true";
defparam \entry_1[49] .power_up = "low";

dffeas \entry_0[49] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[49]~q ),
	.prn(vcc));
defparam \entry_0[49] .is_wysiwyg = "true";
defparam \entry_0[49] .power_up = "low";

dffeas \entry_1[48] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[48]~q ),
	.prn(vcc));
defparam \entry_1[48] .is_wysiwyg = "true";
defparam \entry_1[48] .power_up = "low";

dffeas \entry_0[48] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[48]~q ),
	.prn(vcc));
defparam \entry_0[48] .is_wysiwyg = "true";
defparam \entry_0[48] .power_up = "low";

dffeas \entry_1[51] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[51]~q ),
	.prn(vcc));
defparam \entry_1[51] .is_wysiwyg = "true";
defparam \entry_1[51] .power_up = "low";

dffeas \entry_0[51] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[51]~q ),
	.prn(vcc));
defparam \entry_0[51] .is_wysiwyg = "true";
defparam \entry_0[51] .power_up = "low";

dffeas \entry_1[50] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[50]~q ),
	.prn(vcc));
defparam \entry_1[50] .is_wysiwyg = "true";
defparam \entry_1[50] .power_up = "low";

dffeas \entry_0[50] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[50]~q ),
	.prn(vcc));
defparam \entry_0[50] .is_wysiwyg = "true";
defparam \entry_0[50] .power_up = "low";

dffeas \entry_1[53] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[53]~q ),
	.prn(vcc));
defparam \entry_1[53] .is_wysiwyg = "true";
defparam \entry_1[53] .power_up = "low";

dffeas \entry_0[53] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[53]~q ),
	.prn(vcc));
defparam \entry_0[53] .is_wysiwyg = "true";
defparam \entry_0[53] .power_up = "low";

dffeas \entry_1[52] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[52]~q ),
	.prn(vcc));
defparam \entry_1[52] .is_wysiwyg = "true";
defparam \entry_1[52] .power_up = "low";

dffeas \entry_0[52] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[52]~q ),
	.prn(vcc));
defparam \entry_0[52] .is_wysiwyg = "true";
defparam \entry_0[52] .power_up = "low";

dffeas \entry_1[55] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[55]~q ),
	.prn(vcc));
defparam \entry_1[55] .is_wysiwyg = "true";
defparam \entry_1[55] .power_up = "low";

dffeas \entry_0[55] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[55]~q ),
	.prn(vcc));
defparam \entry_0[55] .is_wysiwyg = "true";
defparam \entry_0[55] .power_up = "low";

dffeas \entry_1[54] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[54]~q ),
	.prn(vcc));
defparam \entry_1[54] .is_wysiwyg = "true";
defparam \entry_1[54] .power_up = "low";

dffeas \entry_0[54] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[54]~q ),
	.prn(vcc));
defparam \entry_0[54] .is_wysiwyg = "true";
defparam \entry_0[54] .power_up = "low";

dffeas \entry_1[57] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[57]~q ),
	.prn(vcc));
defparam \entry_1[57] .is_wysiwyg = "true";
defparam \entry_1[57] .power_up = "low";

dffeas \entry_0[57] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[57]~q ),
	.prn(vcc));
defparam \entry_0[57] .is_wysiwyg = "true";
defparam \entry_0[57] .power_up = "low";

dffeas \entry_1[56] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[56]~q ),
	.prn(vcc));
defparam \entry_1[56] .is_wysiwyg = "true";
defparam \entry_1[56] .power_up = "low";

dffeas \entry_0[56] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[56]~q ),
	.prn(vcc));
defparam \entry_0[56] .is_wysiwyg = "true";
defparam \entry_0[56] .power_up = "low";

dffeas \entry_1[59] (
	.clk(clk),
	.d(src_data_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[59]~q ),
	.prn(vcc));
defparam \entry_1[59] .is_wysiwyg = "true";
defparam \entry_1[59] .power_up = "low";

dffeas \entry_0[59] (
	.clk(clk),
	.d(src_data_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[59]~q ),
	.prn(vcc));
defparam \entry_0[59] .is_wysiwyg = "true";
defparam \entry_0[59] .power_up = "low";

dffeas \entry_1[58] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[58]~q ),
	.prn(vcc));
defparam \entry_1[58] .is_wysiwyg = "true";
defparam \entry_1[58] .power_up = "low";

dffeas \entry_0[58] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[58]~q ),
	.prn(vcc));
defparam \entry_0[58] .is_wysiwyg = "true";
defparam \entry_0[58] .power_up = "low";

dffeas \entry_1[36] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[36]~q ),
	.prn(vcc));
defparam \entry_1[36] .is_wysiwyg = "true";
defparam \entry_1[36] .power_up = "low";

dffeas \entry_0[36] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[36]~q ),
	.prn(vcc));
defparam \entry_0[36] .is_wysiwyg = "true";
defparam \entry_0[36] .power_up = "low";

dffeas \entry_1[37] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[37]~q ),
	.prn(vcc));
defparam \entry_1[37] .is_wysiwyg = "true";
defparam \entry_1[37] .power_up = "low";

dffeas \entry_0[37] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[37]~q ),
	.prn(vcc));
defparam \entry_0[37] .is_wysiwyg = "true";
defparam \entry_0[37] .power_up = "low";

dffeas \entry_1[38] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[38]~q ),
	.prn(vcc));
defparam \entry_1[38] .is_wysiwyg = "true";
defparam \entry_1[38] .power_up = "low";

dffeas \entry_0[38] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[38]~q ),
	.prn(vcc));
defparam \entry_0[38] .is_wysiwyg = "true";
defparam \entry_0[38] .power_up = "low";

dffeas \entry_1[39] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[39]~q ),
	.prn(vcc));
defparam \entry_1[39] .is_wysiwyg = "true";
defparam \entry_1[39] .power_up = "low";

dffeas \entry_0[39] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[39]~q ),
	.prn(vcc));
defparam \entry_0[39] .is_wysiwyg = "true";
defparam \entry_0[39] .power_up = "low";

dffeas \entry_1[40] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[40]~q ),
	.prn(vcc));
defparam \entry_1[40] .is_wysiwyg = "true";
defparam \entry_1[40] .power_up = "low";

dffeas \entry_0[40] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[40]~q ),
	.prn(vcc));
defparam \entry_0[40] .is_wysiwyg = "true";
defparam \entry_0[40] .power_up = "low";

dffeas \entry_1[41] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[41]~q ),
	.prn(vcc));
defparam \entry_1[41] .is_wysiwyg = "true";
defparam \entry_1[41] .power_up = "low";

dffeas \entry_0[41] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[41]~q ),
	.prn(vcc));
defparam \entry_0[41] .is_wysiwyg = "true";
defparam \entry_0[41] .power_up = "low";

dffeas \entry_1[42] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[42]~q ),
	.prn(vcc));
defparam \entry_1[42] .is_wysiwyg = "true";
defparam \entry_1[42] .power_up = "low";

dffeas \entry_0[42] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[42]~q ),
	.prn(vcc));
defparam \entry_0[42] .is_wysiwyg = "true";
defparam \entry_0[42] .power_up = "low";

dffeas \entry_1[43] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[43]~q ),
	.prn(vcc));
defparam \entry_1[43] .is_wysiwyg = "true";
defparam \entry_1[43] .power_up = "low";

dffeas \entry_0[43] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[43]~q ),
	.prn(vcc));
defparam \entry_0[43] .is_wysiwyg = "true";
defparam \entry_0[43] .power_up = "low";

dffeas \entry_1[44] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[44]~q ),
	.prn(vcc));
defparam \entry_1[44] .is_wysiwyg = "true";
defparam \entry_1[44] .power_up = "low";

dffeas \entry_0[44] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[44]~q ),
	.prn(vcc));
defparam \entry_0[44] .is_wysiwyg = "true";
defparam \entry_0[44] .power_up = "low";

dffeas \entry_1[45] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[45]~q ),
	.prn(vcc));
defparam \entry_1[45] .is_wysiwyg = "true";
defparam \entry_1[45] .power_up = "low";

dffeas \entry_0[45] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[45]~q ),
	.prn(vcc));
defparam \entry_0[45] .is_wysiwyg = "true";
defparam \entry_0[45] .power_up = "low";

dffeas \entry_1[32] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[32]~q ),
	.prn(vcc));
defparam \entry_1[32] .is_wysiwyg = "true";
defparam \entry_1[32] .power_up = "low";

dffeas \entry_0[32] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[32]~q ),
	.prn(vcc));
defparam \entry_0[32] .is_wysiwyg = "true";
defparam \entry_0[32] .power_up = "low";

dffeas \entry_1[33] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[33]~q ),
	.prn(vcc));
defparam \entry_1[33] .is_wysiwyg = "true";
defparam \entry_1[33] .power_up = "low";

dffeas \entry_0[33] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[33]~q ),
	.prn(vcc));
defparam \entry_0[33] .is_wysiwyg = "true";
defparam \entry_0[33] .power_up = "low";

dffeas \entry_1[34] (
	.clk(clk),
	.d(comb2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[34]~q ),
	.prn(vcc));
defparam \entry_1[34] .is_wysiwyg = "true";
defparam \entry_1[34] .power_up = "low";

dffeas \entry_0[34] (
	.clk(clk),
	.d(comb2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[34]~q ),
	.prn(vcc));
defparam \entry_0[34] .is_wysiwyg = "true";
defparam \entry_0[34] .power_up = "low";

dffeas \entry_1[35] (
	.clk(clk),
	.d(comb3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[35]~q ),
	.prn(vcc));
defparam \entry_1[35] .is_wysiwyg = "true";
defparam \entry_1[35] .power_up = "low";

dffeas \entry_0[35] (
	.clk(clk),
	.d(comb3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[35]~q ),
	.prn(vcc));
defparam \entry_0[35] .is_wysiwyg = "true";
defparam \entry_0[35] .power_up = "low";

dffeas \entry_1[0] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[0]~q ),
	.prn(vcc));
defparam \entry_1[0] .is_wysiwyg = "true";
defparam \entry_1[0] .power_up = "low";

dffeas \entry_0[0] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[0]~q ),
	.prn(vcc));
defparam \entry_0[0] .is_wysiwyg = "true";
defparam \entry_0[0] .power_up = "low";

dffeas \entry_1[1] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[1]~q ),
	.prn(vcc));
defparam \entry_1[1] .is_wysiwyg = "true";
defparam \entry_1[1] .power_up = "low";

dffeas \entry_0[1] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[1]~q ),
	.prn(vcc));
defparam \entry_0[1] .is_wysiwyg = "true";
defparam \entry_0[1] .power_up = "low";

dffeas \entry_1[2] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[2]~q ),
	.prn(vcc));
defparam \entry_1[2] .is_wysiwyg = "true";
defparam \entry_1[2] .power_up = "low";

dffeas \entry_0[2] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[2]~q ),
	.prn(vcc));
defparam \entry_0[2] .is_wysiwyg = "true";
defparam \entry_0[2] .power_up = "low";

dffeas \entry_1[3] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[3]~q ),
	.prn(vcc));
defparam \entry_1[3] .is_wysiwyg = "true";
defparam \entry_1[3] .power_up = "low";

dffeas \entry_0[3] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[3]~q ),
	.prn(vcc));
defparam \entry_0[3] .is_wysiwyg = "true";
defparam \entry_0[3] .power_up = "low";

dffeas \entry_1[4] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[4]~q ),
	.prn(vcc));
defparam \entry_1[4] .is_wysiwyg = "true";
defparam \entry_1[4] .power_up = "low";

dffeas \entry_0[4] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[4]~q ),
	.prn(vcc));
defparam \entry_0[4] .is_wysiwyg = "true";
defparam \entry_0[4] .power_up = "low";

dffeas \entry_1[5] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[5]~q ),
	.prn(vcc));
defparam \entry_1[5] .is_wysiwyg = "true";
defparam \entry_1[5] .power_up = "low";

dffeas \entry_0[5] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[5]~q ),
	.prn(vcc));
defparam \entry_0[5] .is_wysiwyg = "true";
defparam \entry_0[5] .power_up = "low";

dffeas \entry_1[6] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[6]~q ),
	.prn(vcc));
defparam \entry_1[6] .is_wysiwyg = "true";
defparam \entry_1[6] .power_up = "low";

dffeas \entry_0[6] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[6]~q ),
	.prn(vcc));
defparam \entry_0[6] .is_wysiwyg = "true";
defparam \entry_0[6] .power_up = "low";

dffeas \entry_1[7] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[7]~q ),
	.prn(vcc));
defparam \entry_1[7] .is_wysiwyg = "true";
defparam \entry_1[7] .power_up = "low";

dffeas \entry_0[7] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[7]~q ),
	.prn(vcc));
defparam \entry_0[7] .is_wysiwyg = "true";
defparam \entry_0[7] .power_up = "low";

dffeas \entry_1[8] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[8]~q ),
	.prn(vcc));
defparam \entry_1[8] .is_wysiwyg = "true";
defparam \entry_1[8] .power_up = "low";

dffeas \entry_0[8] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[8]~q ),
	.prn(vcc));
defparam \entry_0[8] .is_wysiwyg = "true";
defparam \entry_0[8] .power_up = "low";

dffeas \entry_1[9] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[9]~q ),
	.prn(vcc));
defparam \entry_1[9] .is_wysiwyg = "true";
defparam \entry_1[9] .power_up = "low";

dffeas \entry_0[9] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[9]~q ),
	.prn(vcc));
defparam \entry_0[9] .is_wysiwyg = "true";
defparam \entry_0[9] .power_up = "low";

dffeas \entry_1[10] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[10]~q ),
	.prn(vcc));
defparam \entry_1[10] .is_wysiwyg = "true";
defparam \entry_1[10] .power_up = "low";

dffeas \entry_0[10] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[10]~q ),
	.prn(vcc));
defparam \entry_0[10] .is_wysiwyg = "true";
defparam \entry_0[10] .power_up = "low";

dffeas \entry_1[11] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[11]~q ),
	.prn(vcc));
defparam \entry_1[11] .is_wysiwyg = "true";
defparam \entry_1[11] .power_up = "low";

dffeas \entry_0[11] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[11]~q ),
	.prn(vcc));
defparam \entry_0[11] .is_wysiwyg = "true";
defparam \entry_0[11] .power_up = "low";

dffeas \entry_1[12] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[12]~q ),
	.prn(vcc));
defparam \entry_1[12] .is_wysiwyg = "true";
defparam \entry_1[12] .power_up = "low";

dffeas \entry_0[12] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[12]~q ),
	.prn(vcc));
defparam \entry_0[12] .is_wysiwyg = "true";
defparam \entry_0[12] .power_up = "low";

dffeas \entry_1[13] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[13]~q ),
	.prn(vcc));
defparam \entry_1[13] .is_wysiwyg = "true";
defparam \entry_1[13] .power_up = "low";

dffeas \entry_0[13] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[13]~q ),
	.prn(vcc));
defparam \entry_0[13] .is_wysiwyg = "true";
defparam \entry_0[13] .power_up = "low";

dffeas \entry_1[14] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[14]~q ),
	.prn(vcc));
defparam \entry_1[14] .is_wysiwyg = "true";
defparam \entry_1[14] .power_up = "low";

dffeas \entry_0[14] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[14]~q ),
	.prn(vcc));
defparam \entry_0[14] .is_wysiwyg = "true";
defparam \entry_0[14] .power_up = "low";

dffeas \entry_1[15] (
	.clk(clk),
	.d(src_payload16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[15]~q ),
	.prn(vcc));
defparam \entry_1[15] .is_wysiwyg = "true";
defparam \entry_1[15] .power_up = "low";

dffeas \entry_0[15] (
	.clk(clk),
	.d(src_payload16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[15]~q ),
	.prn(vcc));
defparam \entry_0[15] .is_wysiwyg = "true";
defparam \entry_0[15] .power_up = "low";

dffeas \entry_1[16] (
	.clk(clk),
	.d(src_payload17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[16]~q ),
	.prn(vcc));
defparam \entry_1[16] .is_wysiwyg = "true";
defparam \entry_1[16] .power_up = "low";

dffeas \entry_0[16] (
	.clk(clk),
	.d(src_payload17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[16]~q ),
	.prn(vcc));
defparam \entry_0[16] .is_wysiwyg = "true";
defparam \entry_0[16] .power_up = "low";

dffeas \entry_1[17] (
	.clk(clk),
	.d(src_payload18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[17]~q ),
	.prn(vcc));
defparam \entry_1[17] .is_wysiwyg = "true";
defparam \entry_1[17] .power_up = "low";

dffeas \entry_0[17] (
	.clk(clk),
	.d(src_payload18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[17]~q ),
	.prn(vcc));
defparam \entry_0[17] .is_wysiwyg = "true";
defparam \entry_0[17] .power_up = "low";

dffeas \entry_1[18] (
	.clk(clk),
	.d(src_payload19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[18]~q ),
	.prn(vcc));
defparam \entry_1[18] .is_wysiwyg = "true";
defparam \entry_1[18] .power_up = "low";

dffeas \entry_0[18] (
	.clk(clk),
	.d(src_payload19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[18]~q ),
	.prn(vcc));
defparam \entry_0[18] .is_wysiwyg = "true";
defparam \entry_0[18] .power_up = "low";

dffeas \entry_1[19] (
	.clk(clk),
	.d(src_payload20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[19]~q ),
	.prn(vcc));
defparam \entry_1[19] .is_wysiwyg = "true";
defparam \entry_1[19] .power_up = "low";

dffeas \entry_0[19] (
	.clk(clk),
	.d(src_payload20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[19]~q ),
	.prn(vcc));
defparam \entry_0[19] .is_wysiwyg = "true";
defparam \entry_0[19] .power_up = "low";

dffeas \entry_1[20] (
	.clk(clk),
	.d(src_payload21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[20]~q ),
	.prn(vcc));
defparam \entry_1[20] .is_wysiwyg = "true";
defparam \entry_1[20] .power_up = "low";

dffeas \entry_0[20] (
	.clk(clk),
	.d(src_payload21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[20]~q ),
	.prn(vcc));
defparam \entry_0[20] .is_wysiwyg = "true";
defparam \entry_0[20] .power_up = "low";

dffeas \entry_1[21] (
	.clk(clk),
	.d(src_payload22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[21]~q ),
	.prn(vcc));
defparam \entry_1[21] .is_wysiwyg = "true";
defparam \entry_1[21] .power_up = "low";

dffeas \entry_0[21] (
	.clk(clk),
	.d(src_payload22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[21]~q ),
	.prn(vcc));
defparam \entry_0[21] .is_wysiwyg = "true";
defparam \entry_0[21] .power_up = "low";

dffeas \entry_1[22] (
	.clk(clk),
	.d(src_payload23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[22]~q ),
	.prn(vcc));
defparam \entry_1[22] .is_wysiwyg = "true";
defparam \entry_1[22] .power_up = "low";

dffeas \entry_0[22] (
	.clk(clk),
	.d(src_payload23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[22]~q ),
	.prn(vcc));
defparam \entry_0[22] .is_wysiwyg = "true";
defparam \entry_0[22] .power_up = "low";

dffeas \entry_1[23] (
	.clk(clk),
	.d(src_payload24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[23]~q ),
	.prn(vcc));
defparam \entry_1[23] .is_wysiwyg = "true";
defparam \entry_1[23] .power_up = "low";

dffeas \entry_0[23] (
	.clk(clk),
	.d(src_payload24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[23]~q ),
	.prn(vcc));
defparam \entry_0[23] .is_wysiwyg = "true";
defparam \entry_0[23] .power_up = "low";

dffeas \entry_1[24] (
	.clk(clk),
	.d(src_payload25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[24]~q ),
	.prn(vcc));
defparam \entry_1[24] .is_wysiwyg = "true";
defparam \entry_1[24] .power_up = "low";

dffeas \entry_0[24] (
	.clk(clk),
	.d(src_payload25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[24]~q ),
	.prn(vcc));
defparam \entry_0[24] .is_wysiwyg = "true";
defparam \entry_0[24] .power_up = "low";

dffeas \entry_1[25] (
	.clk(clk),
	.d(src_payload26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[25]~q ),
	.prn(vcc));
defparam \entry_1[25] .is_wysiwyg = "true";
defparam \entry_1[25] .power_up = "low";

dffeas \entry_0[25] (
	.clk(clk),
	.d(src_payload26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[25]~q ),
	.prn(vcc));
defparam \entry_0[25] .is_wysiwyg = "true";
defparam \entry_0[25] .power_up = "low";

dffeas \entry_1[26] (
	.clk(clk),
	.d(src_payload27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[26]~q ),
	.prn(vcc));
defparam \entry_1[26] .is_wysiwyg = "true";
defparam \entry_1[26] .power_up = "low";

dffeas \entry_0[26] (
	.clk(clk),
	.d(src_payload27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[26]~q ),
	.prn(vcc));
defparam \entry_0[26] .is_wysiwyg = "true";
defparam \entry_0[26] .power_up = "low";

dffeas \entry_1[27] (
	.clk(clk),
	.d(src_payload28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[27]~q ),
	.prn(vcc));
defparam \entry_1[27] .is_wysiwyg = "true";
defparam \entry_1[27] .power_up = "low";

dffeas \entry_0[27] (
	.clk(clk),
	.d(src_payload28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[27]~q ),
	.prn(vcc));
defparam \entry_0[27] .is_wysiwyg = "true";
defparam \entry_0[27] .power_up = "low";

dffeas \entry_1[28] (
	.clk(clk),
	.d(src_payload29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[28]~q ),
	.prn(vcc));
defparam \entry_1[28] .is_wysiwyg = "true";
defparam \entry_1[28] .power_up = "low";

dffeas \entry_0[28] (
	.clk(clk),
	.d(src_payload29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[28]~q ),
	.prn(vcc));
defparam \entry_0[28] .is_wysiwyg = "true";
defparam \entry_0[28] .power_up = "low";

dffeas \entry_1[29] (
	.clk(clk),
	.d(src_payload30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[29]~q ),
	.prn(vcc));
defparam \entry_1[29] .is_wysiwyg = "true";
defparam \entry_1[29] .power_up = "low";

dffeas \entry_0[29] (
	.clk(clk),
	.d(src_payload30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[29]~q ),
	.prn(vcc));
defparam \entry_0[29] .is_wysiwyg = "true";
defparam \entry_0[29] .power_up = "low";

dffeas \entry_1[30] (
	.clk(clk),
	.d(src_payload31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[30]~q ),
	.prn(vcc));
defparam \entry_1[30] .is_wysiwyg = "true";
defparam \entry_1[30] .power_up = "low";

dffeas \entry_0[30] (
	.clk(clk),
	.d(src_payload31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[30]~q ),
	.prn(vcc));
defparam \entry_0[30] .is_wysiwyg = "true";
defparam \entry_0[30] .power_up = "low";

dffeas \entry_1[31] (
	.clk(clk),
	.d(src_payload32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[31]~q ),
	.prn(vcc));
defparam \entry_1[31] .is_wysiwyg = "true";
defparam \entry_1[31] .power_up = "low";

dffeas \entry_0[31] (
	.clk(clk),
	.d(src_payload32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[31]~q ),
	.prn(vcc));
defparam \entry_0[31] .is_wysiwyg = "true";
defparam \entry_0[31] .power_up = "low";

endmodule
