// final_project_soc.v

// Generated using ACDS version 14.1 190 at 2015.05.02.17:56:21

`timescale 1 ps / 1 ps
module final_project_soc (
		inout  wire        audio_config_wire_SDAT,                //              audio_config_wire.SDAT
		output wire        audio_config_wire_SCLK,                //                               .SCLK
		input  wire        audio_wire_ADCDAT,                     //                     audio_wire.ADCDAT
		input  wire        audio_wire_ADCLRCK,                    //                               .ADCLRCK
		input  wire        audio_wire_BCLK,                       //                               .BCLK
		output wire        audio_wire_DACDAT,                     //                               .DACDAT
		input  wire        audio_wire_DACLRCK,                    //                               .DACLRCK
		input  wire        clk_clk,                               //                            clk.clk
		output wire [7:0]  ledg_wire_export,                      //                      ledg_wire.export
		output wire [17:0] ledr_wire_export,                      //                      ledr_wire.export
		input  wire        reset_reset_n,                         //                          reset.reset_n
		output wire        sdram_clk_clk,                         //                      sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                       //                     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                         //                               .ba
		output wire        sdram_wire_cas_n,                      //                               .cas_n
		output wire        sdram_wire_cke,                        //                               .cke
		output wire        sdram_wire_cs_n,                       //                               .cs_n
		inout  wire [31:0] sdram_wire_dq,                         //                               .dq
		output wire [3:0]  sdram_wire_dqm,                        //                               .dqm
		output wire        sdram_wire_ras_n,                      //                               .ras_n
		output wire        sdram_wire_we_n,                       //                               .we_n
		input  wire        unused_sdram_areset_conduit_export,    //    unused_sdram_areset_conduit.export
		output wire        unused_sdram_locked_conduit_export,    //    unused_sdram_locked_conduit.export
		output wire        unused_sdram_phasedone_conduit_export  // unused_sdram_phasedone_conduit.export
	);

	wire         audio_pll_0_audio_clk_clk;                                         // audio_pll_0:audio_clk_clk -> [audio:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:audio_pll_0_audio_clk_clk, rst_controller_001:clk]
	wire         sdram_pll_c0_clk;                                                  // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                 // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                              // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                              // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [28:0] nios2_qsys_0_data_master_address;                                  // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                               // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                     // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                                    // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                          // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                       // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                           // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                              // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;             // mm_interconnect_0:audio_avalon_audio_slave_chipselect -> audio:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;               // audio:readdata -> mm_interconnect_0:audio_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;                // mm_interconnect_0:audio_avalon_audio_slave_address -> audio:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                   // mm_interconnect_0:audio_avalon_audio_slave_read -> audio:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                  // mm_interconnect_0:audio_avalon_audio_slave_write -> audio:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;              // mm_interconnect_0:audio_avalon_audio_slave_writedata -> audio:writedata
	wire  [31:0] mm_interconnect_0_audio_config_avalon_av_config_slave_readdata;    // audio_config:readdata -> mm_interconnect_0:audio_config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_config_avalon_av_config_slave_waitrequest; // audio_config:waitrequest -> mm_interconnect_0:audio_config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_config_avalon_av_config_slave_address;     // mm_interconnect_0:audio_config_avalon_av_config_slave_address -> audio_config:address
	wire         mm_interconnect_0_audio_config_avalon_av_config_slave_read;        // mm_interconnect_0:audio_config_avalon_av_config_slave_read -> audio_config:read
	wire   [3:0] mm_interconnect_0_audio_config_avalon_av_config_slave_byteenable;  // mm_interconnect_0:audio_config_avalon_av_config_slave_byteenable -> audio_config:byteenable
	wire         mm_interconnect_0_audio_config_avalon_av_config_slave_write;       // mm_interconnect_0:audio_config_avalon_av_config_slave_write -> audio_config:write
	wire  [31:0] mm_interconnect_0_audio_config_avalon_av_config_slave_writedata;   // mm_interconnect_0:audio_config_avalon_av_config_slave_writedata -> audio_config:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;          // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;       // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;             // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;              // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;           // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;        // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;            // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;               // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;              // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;          // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;                    // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;                     // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                        // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                       // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;                   // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                             // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                               // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                            // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                   // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                             // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                          // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                  // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                              // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_ledr_s1_chipselect;                              // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                                // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                                 // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                                   // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                               // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                              // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                                // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                                 // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                                   // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                               // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                  // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                    // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;                     // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                  // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                       // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                   // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                       // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver1_irq;                                          // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                              // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         irq_mapper_receiver0_irq;                                          // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                     // audio:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [LEDG:reset_n, LEDR:reset_n, audio_config:reset, audio_pll_0:ref_reset_reset, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [audio:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset]
	wire         audio_pll_0_reset_source_reset;                                    // audio_pll_0:reset_source_reset -> rst_controller_001:reset_in0
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	final_project_soc_LEDG ledg (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_wire_export)                      // external_connection.export
	);

	final_project_soc_LEDR ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_wire_export)                      // external_connection.export
	);

	final_project_soc_audio audio (
		.clk         (audio_pll_0_audio_clk_clk),                             //                clk.clk
		.reset       (rst_controller_001_reset_out_reset),                    //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_synchronizer_receiver_irq),                         //          interrupt.irq
		.AUD_ADCDAT  (audio_wire_ADCDAT),                                     // external_interface.export
		.AUD_ADCLRCK (audio_wire_ADCLRCK),                                    //                   .export
		.AUD_BCLK    (audio_wire_BCLK),                                       //                   .export
		.AUD_DACDAT  (audio_wire_DACDAT),                                     //                   .export
		.AUD_DACLRCK (audio_wire_DACLRCK)                                     //                   .export
	);

	final_project_soc_audio_config audio_config (
		.clk         (clk_clk),                                                           //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                    //                  reset.reset
		.address     (mm_interconnect_0_audio_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_config_wire_SDAT),                                            //     external_interface.export
		.I2C_SCLK    (audio_config_wire_SCLK)                                             //                       .export
	);

	final_project_soc_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (rst_controller_reset_out_reset), //    ref_reset.reset
		.audio_clk_clk      (audio_pll_0_audio_clk_clk),      //    audio_clk.clk
		.reset_source_reset (audio_pll_0_reset_source_reset)  // reset_source.reset
	);

	final_project_soc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	final_project_soc_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	final_project_soc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	final_project_soc_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_project_soc_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                   //                    c1.clk
		.areset    (unused_sdram_areset_conduit_export),              //        areset_conduit.export
		.locked    (unused_sdram_locked_conduit_export),              //        locked_conduit.export
		.phasedone (unused_sdram_phasedone_conduit_export)            //     phasedone_conduit.export
	);

	final_project_soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	final_project_soc_mm_interconnect_0 mm_interconnect_0 (
		.audio_pll_0_audio_clk_clk                       (audio_pll_0_audio_clk_clk),                                         //                    audio_pll_0_audio_clk.clk
		.clk_0_clk_clk                                   (clk_clk),                                                           //                                clk_0_clk.clk
		.sdram_pll_c0_clk                                (sdram_pll_c0_clk),                                                  //                             sdram_pll_c0.clk
		.audio_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                                //        audio_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                    // nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset         (rst_controller_002_reset_out_reset),                                //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                (nios2_qsys_0_data_master_address),                                  //                 nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest            (nios2_qsys_0_data_master_waitrequest),                              //                                         .waitrequest
		.nios2_qsys_0_data_master_byteenable             (nios2_qsys_0_data_master_byteenable),                               //                                         .byteenable
		.nios2_qsys_0_data_master_read                   (nios2_qsys_0_data_master_read),                                     //                                         .read
		.nios2_qsys_0_data_master_readdata               (nios2_qsys_0_data_master_readdata),                                 //                                         .readdata
		.nios2_qsys_0_data_master_write                  (nios2_qsys_0_data_master_write),                                    //                                         .write
		.nios2_qsys_0_data_master_writedata              (nios2_qsys_0_data_master_writedata),                                //                                         .writedata
		.nios2_qsys_0_data_master_debugaccess            (nios2_qsys_0_data_master_debugaccess),                              //                                         .debugaccess
		.nios2_qsys_0_instruction_master_address         (nios2_qsys_0_instruction_master_address),                           //          nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest     (nios2_qsys_0_instruction_master_waitrequest),                       //                                         .waitrequest
		.nios2_qsys_0_instruction_master_read            (nios2_qsys_0_instruction_master_read),                              //                                         .read
		.nios2_qsys_0_instruction_master_readdata        (nios2_qsys_0_instruction_master_readdata),                          //                                         .readdata
		.audio_avalon_audio_slave_address                (mm_interconnect_0_audio_avalon_audio_slave_address),                //                 audio_avalon_audio_slave.address
		.audio_avalon_audio_slave_write                  (mm_interconnect_0_audio_avalon_audio_slave_write),                  //                                         .write
		.audio_avalon_audio_slave_read                   (mm_interconnect_0_audio_avalon_audio_slave_read),                   //                                         .read
		.audio_avalon_audio_slave_readdata               (mm_interconnect_0_audio_avalon_audio_slave_readdata),               //                                         .readdata
		.audio_avalon_audio_slave_writedata              (mm_interconnect_0_audio_avalon_audio_slave_writedata),              //                                         .writedata
		.audio_avalon_audio_slave_chipselect             (mm_interconnect_0_audio_avalon_audio_slave_chipselect),             //                                         .chipselect
		.audio_config_avalon_av_config_slave_address     (mm_interconnect_0_audio_config_avalon_av_config_slave_address),     //      audio_config_avalon_av_config_slave.address
		.audio_config_avalon_av_config_slave_write       (mm_interconnect_0_audio_config_avalon_av_config_slave_write),       //                                         .write
		.audio_config_avalon_av_config_slave_read        (mm_interconnect_0_audio_config_avalon_av_config_slave_read),        //                                         .read
		.audio_config_avalon_av_config_slave_readdata    (mm_interconnect_0_audio_config_avalon_av_config_slave_readdata),    //                                         .readdata
		.audio_config_avalon_av_config_slave_writedata   (mm_interconnect_0_audio_config_avalon_av_config_slave_writedata),   //                                         .writedata
		.audio_config_avalon_av_config_slave_byteenable  (mm_interconnect_0_audio_config_avalon_av_config_slave_byteenable),  //                                         .byteenable
		.audio_config_avalon_av_config_slave_waitrequest (mm_interconnect_0_audio_config_avalon_av_config_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),           //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),             //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),              //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),          //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),         //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),       //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),        //                                         .chipselect
		.LEDG_s1_address                                 (mm_interconnect_0_ledg_s1_address),                                 //                                  LEDG_s1.address
		.LEDG_s1_write                                   (mm_interconnect_0_ledg_s1_write),                                   //                                         .write
		.LEDG_s1_readdata                                (mm_interconnect_0_ledg_s1_readdata),                                //                                         .readdata
		.LEDG_s1_writedata                               (mm_interconnect_0_ledg_s1_writedata),                               //                                         .writedata
		.LEDG_s1_chipselect                              (mm_interconnect_0_ledg_s1_chipselect),                              //                                         .chipselect
		.LEDR_s1_address                                 (mm_interconnect_0_ledr_s1_address),                                 //                                  LEDR_s1.address
		.LEDR_s1_write                                   (mm_interconnect_0_ledr_s1_write),                                   //                                         .write
		.LEDR_s1_readdata                                (mm_interconnect_0_ledr_s1_readdata),                                //                                         .readdata
		.LEDR_s1_writedata                               (mm_interconnect_0_ledr_s1_writedata),                               //                                         .writedata
		.LEDR_s1_chipselect                              (mm_interconnect_0_ledr_s1_chipselect),                              //                                         .chipselect
		.nios2_qsys_0_debug_mem_slave_address            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),            //             nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),              //                                         .write
		.nios2_qsys_0_debug_mem_slave_read               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),               //                                         .read
		.nios2_qsys_0_debug_mem_slave_readdata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),           //                                         .readdata
		.nios2_qsys_0_debug_mem_slave_writedata          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),          //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),         //                                         .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest        (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),        //                                         .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess        (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),        //                                         .debugaccess
		.onchip_memory2_0_s1_address                     (mm_interconnect_0_onchip_memory2_0_s1_address),                     //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                       (mm_interconnect_0_onchip_memory2_0_s1_write),                       //                                         .write
		.onchip_memory2_0_s1_readdata                    (mm_interconnect_0_onchip_memory2_0_s1_readdata),                    //                                         .readdata
		.onchip_memory2_0_s1_writedata                   (mm_interconnect_0_onchip_memory2_0_s1_writedata),                   //                                         .writedata
		.onchip_memory2_0_s1_byteenable                  (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                  //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                  (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                  //                                         .chipselect
		.onchip_memory2_0_s1_clken                       (mm_interconnect_0_onchip_memory2_0_s1_clken),                       //                                         .clken
		.sdram_s1_address                                (mm_interconnect_0_sdram_s1_address),                                //                                 sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_0_sdram_s1_write),                                  //                                         .write
		.sdram_s1_read                                   (mm_interconnect_0_sdram_s1_read),                                   //                                         .read
		.sdram_s1_readdata                               (mm_interconnect_0_sdram_s1_readdata),                               //                                         .readdata
		.sdram_s1_writedata                              (mm_interconnect_0_sdram_s1_writedata),                              //                                         .writedata
		.sdram_s1_byteenable                             (mm_interconnect_0_sdram_s1_byteenable),                             //                                         .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_0_sdram_s1_readdatavalid),                          //                                         .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_0_sdram_s1_waitrequest),                            //                                         .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_0_sdram_s1_chipselect),                             //                                         .chipselect
		.sdram_pll_pll_slave_address                     (mm_interconnect_0_sdram_pll_pll_slave_address),                     //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                       (mm_interconnect_0_sdram_pll_pll_slave_write),                       //                                         .write
		.sdram_pll_pll_slave_read                        (mm_interconnect_0_sdram_pll_pll_slave_read),                        //                                         .read
		.sdram_pll_pll_slave_readdata                    (mm_interconnect_0_sdram_pll_pll_slave_readdata),                    //                                         .readdata
		.sdram_pll_pll_slave_writedata                   (mm_interconnect_0_sdram_pll_pll_slave_writedata),                   //                                         .writedata
		.sysid_qsys_0_control_slave_address              (mm_interconnect_0_sysid_qsys_0_control_slave_address),              //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata             (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)              //                                         .readdata
	);

	final_project_soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_0_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (audio_pll_0_audio_clk_clk),          //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (audio_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (audio_pll_0_audio_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
