// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 14.1.1 Build 190 01/19/2015 SJ Web Edition"

// DATE "05/01/2015 22:30:07"

// 
// Device: Altera EP4CE115F29C7 Package FBGA780
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module final_project_soc (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	audio_config_wire_SDAT,
	audio_config_wire_SCLK,
	audio_wire_ADCDAT,
	audio_wire_ADCLRCK,
	audio_wire_BCLK,
	audio_wire_DACDAT,
	audio_wire_DACLRCK,
	clk_clk,
	ledg_wire_export,
	ledr_wire_export,
	reset_reset_n,
	sdram_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	unused_sdram_areset_conduit_export,
	unused_sdram_locked_conduit_export,
	unused_sdram_phasedone_conduit_export)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
inout 	audio_config_wire_SDAT;
output 	audio_config_wire_SCLK;
input 	audio_wire_ADCDAT;
input 	audio_wire_ADCLRCK;
input 	audio_wire_BCLK;
output 	audio_wire_DACDAT;
input 	audio_wire_DACLRCK;
input 	clk_clk;
output 	[7:0] ledg_wire_export;
output 	[17:0] ledr_wire_export;
input 	reset_reset_n;
output 	sdram_clk_clk;
output 	[12:0] sdram_wire_addr;
output 	[1:0] sdram_wire_ba;
output 	sdram_wire_cas_n;
output 	sdram_wire_cke;
output 	sdram_wire_cs_n;
inout 	[31:0] sdram_wire_dq;
output 	[3:0] sdram_wire_dqm;
output 	sdram_wire_ras_n;
output 	sdram_wire_we_n;
input 	unused_sdram_areset_conduit_export;
output 	unused_sdram_locked_conduit_export;
output 	unused_sdram_phasedone_conduit_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdram_pll|sd1|wire_pll7_clk[0] ;
wire \sdram_pll|sd1|wire_pll7_clk[1] ;
wire \sdram|m_addr[0]~q ;
wire \sdram|m_addr[1]~q ;
wire \sdram|m_addr[2]~q ;
wire \sdram|m_addr[3]~q ;
wire \sdram|m_addr[4]~q ;
wire \sdram|m_addr[5]~q ;
wire \sdram|m_addr[6]~q ;
wire \sdram|m_addr[7]~q ;
wire \sdram|m_addr[8]~q ;
wire \sdram|m_addr[9]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[0]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[28]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[27]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[26]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[25]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[24]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[23]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[22]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[21]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[20]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[19]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[18]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[17]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[16]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[15]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[14]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[13]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[6]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[7]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[5]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[4]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[12]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[10]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[9]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[8]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[11]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[2]~q ;
wire \nios2_qsys_0|cpu|W_alu_result[3]~q ;
wire \audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|locked ;
wire \audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|clk[0] ;
wire \sdram|oe~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ;
wire \audio_config|readdata[0]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ;
wire \audio_config|readdata[1]~q ;
wire \audio_config|readdata[2]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ;
wire \audio_config|readdata[16]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ;
wire \audio_config|readdata[17]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ;
wire \audio_config|readdata[8]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[0]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[1]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[2]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[3]~q ;
wire \nios2_qsys_0|cpu|d_writedata[31]~q ;
wire \nios2_qsys_0|cpu|d_writedata[30]~q ;
wire \nios2_qsys_0|cpu|d_writedata[29]~q ;
wire \nios2_qsys_0|cpu|d_writedata[28]~q ;
wire \nios2_qsys_0|cpu|d_writedata[27]~q ;
wire \nios2_qsys_0|cpu|d_writedata[26]~q ;
wire \nios2_qsys_0|cpu|d_writedata[25]~q ;
wire \nios2_qsys_0|cpu|d_writedata[24]~q ;
wire \audio|readdata[0]~q ;
wire \audio|readdata[1]~q ;
wire \audio|readdata[2]~q ;
wire \audio|readdata[3]~q ;
wire \audio|readdata[4]~q ;
wire \audio|readdata[11]~q ;
wire \audio|readdata[13]~q ;
wire \audio|readdata[16]~q ;
wire \audio|readdata[12]~q ;
wire \audio|readdata[5]~q ;
wire \audio|readdata[14]~q ;
wire \audio|readdata[15]~q ;
wire \audio|readdata[21]~q ;
wire \audio|readdata[18]~q ;
wire \audio|readdata[17]~q ;
wire \audio|readdata[31]~q ;
wire \audio|readdata[30]~q ;
wire \audio|readdata[29]~q ;
wire \audio|readdata[28]~q ;
wire \audio|readdata[27]~q ;
wire \audio|readdata[26]~q ;
wire \audio|readdata[25]~q ;
wire \audio|readdata[10]~q ;
wire \audio|readdata[24]~q ;
wire \audio|readdata[9]~q ;
wire \audio|readdata[23]~q ;
wire \audio|readdata[8]~q ;
wire \audio|readdata[22]~q ;
wire \audio|readdata[7]~q ;
wire \audio|readdata[6]~q ;
wire \audio|readdata[20]~q ;
wire \audio|readdata[19]~q ;
wire \audio|irq~q ;
wire \audio_config|Serial_Bus_Controller|serial_clk~0_combout ;
wire \audio|Audio_Out_Serializer|serial_audio_out_data~q ;
wire \ledg|data_out[0]~q ;
wire \ledg|data_out[1]~q ;
wire \ledg|data_out[2]~q ;
wire \ledg|data_out[3]~q ;
wire \ledg|data_out[4]~q ;
wire \ledg|data_out[5]~q ;
wire \ledg|data_out[6]~q ;
wire \ledg|data_out[7]~q ;
wire \ledr|data_out[0]~q ;
wire \ledr|data_out[1]~q ;
wire \ledr|data_out[2]~q ;
wire \ledr|data_out[3]~q ;
wire \ledr|data_out[4]~q ;
wire \ledr|data_out[5]~q ;
wire \ledr|data_out[6]~q ;
wire \ledr|data_out[7]~q ;
wire \ledr|data_out[8]~q ;
wire \ledr|data_out[9]~q ;
wire \ledr|data_out[10]~q ;
wire \ledr|data_out[11]~q ;
wire \ledr|data_out[12]~q ;
wire \ledr|data_out[13]~q ;
wire \ledr|data_out[14]~q ;
wire \ledr|data_out[15]~q ;
wire \ledr|data_out[16]~q ;
wire \ledr|data_out[17]~q ;
wire \sdram|m_addr[10]~q ;
wire \sdram|m_addr[11]~q ;
wire \sdram|m_addr[12]~q ;
wire \sdram|m_bank[0]~q ;
wire \sdram|m_bank[1]~q ;
wire \sdram|m_cmd[1]~q ;
wire \sdram|m_cmd[3]~q ;
wire \sdram|m_dqm[0]~q ;
wire \sdram|m_dqm[1]~q ;
wire \sdram|m_dqm[2]~q ;
wire \sdram|m_dqm[3]~q ;
wire \sdram|m_cmd[2]~q ;
wire \sdram|m_cmd[0]~q ;
wire \sdram_pll|sd1|locked~combout ;
wire \jtag_uart_0|final_project_soc_jtag_uart_0_alt_jtag_atlantic|tdo~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|ir_out[0]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|ir_out[1]~q ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[1]~q ;
wire \nios2_qsys_0|cpu|d_read~q ;
wire \nios2_qsys_0|cpu|d_write~q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_translator|read_accepted~q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_translator|write_accepted~q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_agent|cp_valid~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_valid~1_combout ;
wire \nios2_qsys_0|cpu|F_pc[26]~q ;
wire \nios2_qsys_0|cpu|F_pc[25]~q ;
wire \nios2_qsys_0|cpu|F_pc[24]~q ;
wire \nios2_qsys_0|cpu|F_pc[23]~q ;
wire \nios2_qsys_0|cpu|F_pc[22]~q ;
wire \nios2_qsys_0|cpu|F_pc[21]~q ;
wire \nios2_qsys_0|cpu|F_pc[20]~q ;
wire \nios2_qsys_0|cpu|F_pc[19]~q ;
wire \nios2_qsys_0|cpu|F_pc[18]~q ;
wire \nios2_qsys_0|cpu|F_pc[17]~q ;
wire \nios2_qsys_0|cpu|F_pc[16]~q ;
wire \nios2_qsys_0|cpu|F_pc[15]~q ;
wire \nios2_qsys_0|cpu|F_pc[14]~q ;
wire \nios2_qsys_0|cpu|F_pc[13]~q ;
wire \nios2_qsys_0|cpu|F_pc[12]~q ;
wire \nios2_qsys_0|cpu|F_pc[11]~q ;
wire \nios2_qsys_0|cpu|F_pc[10]~q ;
wire \nios2_qsys_0|cpu|F_pc[8]~q ;
wire \nios2_qsys_0|cpu|F_pc[7]~q ;
wire \nios2_qsys_0|cpu|F_pc[6]~q ;
wire \nios2_qsys_0|cpu|F_pc[5]~q ;
wire \nios2_qsys_0|cpu|F_pc[3]~q ;
wire \nios2_qsys_0|cpu|i_read~q ;
wire \nios2_qsys_0|cpu|F_pc[2]~q ;
wire \nios2_qsys_0|cpu|F_pc[4]~q ;
wire \nios2_qsys_0|cpu|F_pc[9]~q ;
wire \mm_interconnect_0|cmd_demux_001|src1_valid~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_write~0_combout ;
wire \mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \audio_config|internal_reset~2_combout ;
wire \nios2_qsys_0|cpu|d_writedata[0]~q ;
wire \nios2_qsys_0|cpu|d_byteenable[0]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[32]~combout ;
wire \nios2_qsys_0|cpu|F_pc[0]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[38]~combout ;
wire \nios2_qsys_0|cpu|F_pc[1]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[39]~combout ;
wire \rst_controller|r_sync_rst~q ;
wire \rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|router|Equal0~2_combout ;
wire \mm_interconnect_0|ledg_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \ledg|always0~0_combout ;
wire \ledg|always0~1_combout ;
wire \mm_interconnect_0|ledg_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|ledg_s1_translator|wait_latency_counter[0]~q ;
wire \nios2_qsys_0|cpu|d_writedata[1]~q ;
wire \nios2_qsys_0|cpu|d_writedata[2]~q ;
wire \nios2_qsys_0|cpu|d_writedata[3]~q ;
wire \nios2_qsys_0|cpu|d_writedata[4]~q ;
wire \nios2_qsys_0|cpu|d_writedata[5]~q ;
wire \nios2_qsys_0|cpu|d_writedata[6]~q ;
wire \nios2_qsys_0|cpu|d_writedata[7]~q ;
wire \mm_interconnect_0|router|Equal2~1_combout ;
wire \mm_interconnect_0|ledr_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \ledr|always0~0_combout ;
wire \mm_interconnect_0|ledr_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|ledr_s1_translator|wait_latency_counter[0]~q ;
wire \nios2_qsys_0|cpu|d_writedata[8]~q ;
wire \nios2_qsys_0|cpu|d_writedata[9]~q ;
wire \nios2_qsys_0|cpu|d_writedata[10]~q ;
wire \nios2_qsys_0|cpu|d_writedata[11]~q ;
wire \nios2_qsys_0|cpu|d_writedata[12]~q ;
wire \nios2_qsys_0|cpu|d_writedata[13]~q ;
wire \nios2_qsys_0|cpu|d_writedata[14]~q ;
wire \nios2_qsys_0|cpu|d_writedata[15]~q ;
wire \nios2_qsys_0|cpu|d_writedata[16]~q ;
wire \nios2_qsys_0|cpu|d_writedata[17]~q ;
wire \sdram|the_final_project_soc_sdram_input_efifo_module|entries[1]~q ;
wire \sdram|the_final_project_soc_sdram_input_efifo_module|entries[0]~q ;
wire \rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|cmd_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_read~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[68]~combout ;
wire \audio_config|waitrequest~1_combout ;
wire \audio_config|Equal2~0_combout ;
wire \audio_config|s_serial_transfer.STATE_1_PRE_WRITE~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|audio_config_avalon_av_config_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_toggle_flopped~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|ledg_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|ledr_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ;
wire \mm_interconnect_0|sdram_pll_pll_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_009|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|ledr_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[67]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[67]~q ;
wire \mm_interconnect_0|ledg_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~0_combout ;
wire \jtag_uart_0|final_project_soc_jtag_uart_0_alt_jtag_atlantic|rst1~q ;
wire \mm_interconnect_0|router|Equal2~4_combout ;
wire \jtag_uart_0|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_009|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \audio_config|waitrequest~combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_translator|av_waitrequest~2_combout ;
wire \mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_004|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_009|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_valid~combout ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_agent|av_readdatavalid~4_combout ;
wire \mm_interconnect_0|cmd_mux|saved_grant[0]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[3]~q ;
wire \mm_interconnect_0|cmd_mux|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux|WideOr1~combout ;
wire \mm_interconnect_0|audio_avalon_audio_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux|last_cycle~0_combout ;
wire \mm_interconnect_0|audio_avalon_audio_slave_agent|nonposted_write_endofpacket~0_combout ;
wire \mm_interconnect_0|cmd_mux_005|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[38]~combout ;
wire \mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem~0_combout ;
wire \mm_interconnect_0|cmd_mux_005|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_006|last_cycle~0_combout ;
wire \mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ;
wire \mm_interconnect_0|cmd_mux_006|WideOr1~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[68]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[62]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[51]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[50]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[53]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[52]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[55]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[54]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[57]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[56]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[59]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[58]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[61]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[60]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_006|src_data[47]~combout ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[32]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[32]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[33]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[33]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[34]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[34]~q ;
wire \mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[35]~q ;
wire \mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[35]~q ;
wire \audio_config|Serial_Bus_Controller|serial_data~1_combout ;
wire \audio_config|Serial_Bus_Controller|serial_data~2_combout ;
wire \sdram|m_data[0]~q ;
wire \sdram|m_data[1]~q ;
wire \sdram|m_data[2]~q ;
wire \sdram|m_data[3]~q ;
wire \sdram|m_data[4]~q ;
wire \sdram|m_data[5]~q ;
wire \sdram|m_data[6]~q ;
wire \sdram|m_data[7]~q ;
wire \sdram|m_data[8]~q ;
wire \sdram|m_data[9]~q ;
wire \sdram|m_data[10]~q ;
wire \sdram|m_data[11]~q ;
wire \sdram|m_data[12]~q ;
wire \sdram|m_data[13]~q ;
wire \sdram|m_data[14]~q ;
wire \sdram|m_data[15]~q ;
wire \sdram|m_data[16]~q ;
wire \sdram|m_data[17]~q ;
wire \sdram|m_data[18]~q ;
wire \sdram|m_data[19]~q ;
wire \sdram|m_data[20]~q ;
wire \sdram|m_data[21]~q ;
wire \sdram|m_data[22]~q ;
wire \sdram|m_data[23]~q ;
wire \sdram|m_data[24]~q ;
wire \sdram|m_data[25]~q ;
wire \sdram|m_data[26]~q ;
wire \sdram|m_data[27]~q ;
wire \sdram|m_data[28]~q ;
wire \sdram|m_data[29]~q ;
wire \sdram|m_data[30]~q ;
wire \sdram|m_data[31]~q ;
wire \mm_interconnect_0|audio_config_avalon_av_config_slave_agent|m0_read~combout ;
wire \mm_interconnect_0|cmd_mux_004|WideOr1~combout ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent|local_read~0_combout ;
wire \mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem~1_combout ;
wire \mm_interconnect_0|cmd_mux_009|WideOr1~combout ;
wire \nios2_qsys_0|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|sdram_pll_pll_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[0]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[0]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[1]~q ;
wire \mm_interconnect_0|sdram_pll_pll_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[1]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[2]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[2]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \audio_config|readdata[3]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[3]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[3]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \audio_config|readdata[4]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[4]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[4]~q ;
wire \mm_interconnect_0|cmd_mux|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux|src_data[68]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~0_combout ;
wire \nios2_qsys_0|cpu|d_byteenable[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem~4_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[46]~combout ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[11]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[11]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[13]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[13]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~3_combout ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[16]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[16]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[12]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[12]~q ;
wire \audio_config|readdata[5]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[5]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[5]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[14]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[14]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[15]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[15]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[21]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[21]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[18]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[18]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[17]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[17]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[31]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[31]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[28]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[28]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[27]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[27]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[26]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[26]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[10]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[10]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[24]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[24]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[9]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[9]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[23]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[23]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[8]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[8]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[22]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[22]~q ;
wire \audio_config|readdata[7]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[7]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[7]~q ;
wire \audio_config|readdata[6]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[6]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[6]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[20]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[20]~q ;
wire \mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[19]~q ;
wire \mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[19]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~9_combout ;
wire \jtag_uart_0|av_readdata[9]~combout ;
wire \jtag_uart_0|av_readdata[8]~0_combout ;
wire \irq_synchronizer|sync|sync[0].u|dreg[1]~q ;
wire \rst_controller|r_early_rst~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[32]~combout ;
wire \sdram_pll|readdata[0]~1_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~1_combout ;
wire \sdram_pll|readdata[1]~2_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~3_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[4]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~11_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~14_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~16_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~19_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~21_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~24_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~26_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~29_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~32_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~35_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~38_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~41_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[10]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[16]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[17]~combout ;
wire \nios2_qsys_0|cpu|d_byteenable[1]~q ;
wire \nios2_qsys_0|cpu|d_byteenable[3]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_006|src_payload~32_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[11]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[33]~combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[13]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[34]~combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[16]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~8_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[12]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~9_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[5]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~10_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[14]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[15]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~11_combout ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[28]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[28]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[21]~q ;
wire \nios2_qsys_0|cpu|d_writedata[21]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~12_combout ;
wire \nios2_qsys_0|cpu|d_writedata[18]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~13_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[18]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[27]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[27]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[17]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_data[35]~combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[31]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[26]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[26]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~16_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[30]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[25]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~17_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[29]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[24]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[24]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~18_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[28]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[23]~73_combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~19_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[27]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[22]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~20_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[26]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[21]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~21_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[25]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[20]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~22_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[10]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~23_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[24]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[19]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~24_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[9]~q ;
wire \nios2_qsys_0|cpu|d_writedata[23]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~25_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[23]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[18]~combout ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~26_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[8]~q ;
wire \nios2_qsys_0|cpu|d_writedata[22]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~27_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[22]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~28_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[7]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~29_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[6]~q ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[20]~q ;
wire \nios2_qsys_0|cpu|d_writedata[20]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~30_combout ;
wire \nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[19]~q ;
wire \nios2_qsys_0|cpu|d_writedata[19]~q ;
wire \mm_interconnect_0|cmd_mux_009|src_payload~31_combout ;
wire \ledr|readdata[0]~combout ;
wire \jtag_uart_0|read_0~q ;
wire \jtag_uart_0|av_readdata[0]~1_combout ;
wire \ledg|readdata[0]~combout ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \mm_interconnect_0|cmd_mux|src_payload~2_combout ;
wire \ledr|readdata[1]~combout ;
wire \jtag_uart_0|av_readdata[1]~2_combout ;
wire \ledg|readdata[1]~combout ;
wire \ledr|readdata[2]~combout ;
wire \jtag_uart_0|av_readdata[2]~3_combout ;
wire \ledg|readdata[2]~combout ;
wire \ledr|readdata[3]~combout ;
wire \jtag_uart_0|av_readdata[3]~4_combout ;
wire \ledg|readdata[3]~combout ;
wire \ledr|readdata[4]~combout ;
wire \jtag_uart_0|av_readdata[4]~5_combout ;
wire \ledg|readdata[4]~combout ;
wire \ledr|readdata[5]~combout ;
wire \jtag_uart_0|av_readdata[5]~6_combout ;
wire \ledg|readdata[5]~combout ;
wire \ledr|readdata[6]~combout ;
wire \jtag_uart_0|av_readdata[6]~7_combout ;
wire \ledg|readdata[6]~combout ;
wire \ledr|readdata[7]~combout ;
wire \jtag_uart_0|av_readdata[7]~8_combout ;
wire \ledg|readdata[7]~combout ;
wire \ledr|readdata[8]~combout ;
wire \ledr|readdata[9]~combout ;
wire \ledr|readdata[10]~combout ;
wire \jtag_uart_0|ac~q ;
wire \ledr|readdata[11]~combout ;
wire \ledr|readdata[12]~combout ;
wire \ledr|readdata[13]~combout ;
wire \ledr|readdata[14]~combout ;
wire \jtag_uart_0|woverflow~q ;
wire \ledr|readdata[15]~combout ;
wire \jtag_uart_0|rvalid~q ;
wire \ledr|readdata[16]~combout ;
wire \ledr|readdata[17]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[32]~combout ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[31]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[31]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[30]~q ;
wire \mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[29]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~3_combout ;
wire \sdram|za_valid~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[0]~q ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[1]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~4_combout ;
wire \mm_interconnect_0|crosser|clock_xer|out_data_buffer[2]~q ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_004|src_payload~32_combout ;
wire \sdram|za_data[0]~q ;
wire \sdram|za_data[1]~q ;
wire \sdram|za_data[2]~q ;
wire \sdram|za_data[3]~q ;
wire \sdram|za_data[4]~q ;
wire \mm_interconnect_0|cmd_mux|src_payload~5_combout ;
wire \sdram|za_data[11]~q ;
wire \sdram|za_data[13]~q ;
wire \sdram|za_data[16]~q ;
wire \sdram|za_data[12]~q ;
wire \sdram|za_data[5]~q ;
wire \sdram|za_data[14]~q ;
wire \sdram|za_data[15]~q ;
wire \sdram|za_data[21]~q ;
wire \sdram|za_data[18]~q ;
wire \sdram|za_data[17]~q ;
wire \sdram|za_data[31]~q ;
wire \sdram|za_data[30]~q ;
wire \sdram|za_data[29]~q ;
wire \sdram|za_data[28]~q ;
wire \sdram|za_data[27]~q ;
wire \sdram|za_data[26]~q ;
wire \sdram|za_data[25]~q ;
wire \sdram|za_data[10]~q ;
wire \sdram|za_data[24]~q ;
wire \sdram|za_data[9]~q ;
wire \sdram|za_data[23]~q ;
wire \sdram|za_data[8]~q ;
wire \sdram|za_data[22]~q ;
wire \sdram|za_data[7]~q ;
wire \sdram|za_data[6]~q ;
wire \sdram|za_data[20]~q ;
wire \sdram|za_data[19]~q ;
wire \mm_interconnect_0|cmd_mux|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux|src_payload~31_combout ;
wire \nios2_qsys_0|cpu|av_ld_getting_data~9_combout ;
wire \mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~84_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~85_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \audio_config_wire_SDAT~input_o ;
wire \sdram_wire_dq[0]~input_o ;
wire \sdram_wire_dq[1]~input_o ;
wire \sdram_wire_dq[2]~input_o ;
wire \sdram_wire_dq[3]~input_o ;
wire \sdram_wire_dq[4]~input_o ;
wire \sdram_wire_dq[5]~input_o ;
wire \sdram_wire_dq[6]~input_o ;
wire \sdram_wire_dq[7]~input_o ;
wire \sdram_wire_dq[8]~input_o ;
wire \sdram_wire_dq[9]~input_o ;
wire \sdram_wire_dq[10]~input_o ;
wire \sdram_wire_dq[11]~input_o ;
wire \sdram_wire_dq[12]~input_o ;
wire \sdram_wire_dq[13]~input_o ;
wire \sdram_wire_dq[14]~input_o ;
wire \sdram_wire_dq[15]~input_o ;
wire \sdram_wire_dq[16]~input_o ;
wire \sdram_wire_dq[17]~input_o ;
wire \sdram_wire_dq[18]~input_o ;
wire \sdram_wire_dq[19]~input_o ;
wire \sdram_wire_dq[20]~input_o ;
wire \sdram_wire_dq[21]~input_o ;
wire \sdram_wire_dq[22]~input_o ;
wire \sdram_wire_dq[23]~input_o ;
wire \sdram_wire_dq[24]~input_o ;
wire \sdram_wire_dq[25]~input_o ;
wire \sdram_wire_dq[26]~input_o ;
wire \sdram_wire_dq[27]~input_o ;
wire \sdram_wire_dq[28]~input_o ;
wire \sdram_wire_dq[29]~input_o ;
wire \sdram_wire_dq[30]~input_o ;
wire \sdram_wire_dq[31]~input_o ;
wire \clk_clk~input_o ;
wire \unused_sdram_areset_conduit_export~input_o ;
wire \reset_reset_n~input_o ;
wire \audio_wire_DACLRCK~input_o ;
wire \audio_wire_BCLK~input_o ;
wire \audio_wire_ADCLRCK~input_o ;
wire \audio_wire_ADCDAT~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;


final_project_soc_final_project_soc_LEDR ledr(
	.W_alu_result_6(\nios2_qsys_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_2(\nios2_qsys_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_qsys_0|cpu|W_alu_result[3]~q ),
	.data_out_0(\ledr|data_out[0]~q ),
	.data_out_1(\ledr|data_out[1]~q ),
	.data_out_2(\ledr|data_out[2]~q ),
	.data_out_3(\ledr|data_out[3]~q ),
	.data_out_4(\ledr|data_out[4]~q ),
	.data_out_5(\ledr|data_out[5]~q ),
	.data_out_6(\ledr|data_out[6]~q ),
	.data_out_7(\ledr|data_out[7]~q ),
	.data_out_8(\ledr|data_out[8]~q ),
	.data_out_9(\ledr|data_out[9]~q ),
	.data_out_10(\ledr|data_out[10]~q ),
	.data_out_11(\ledr|data_out[11]~q ),
	.data_out_12(\ledr|data_out[12]~q ),
	.data_out_13(\ledr|data_out[13]~q ),
	.data_out_14(\ledr|data_out[14]~q ),
	.data_out_15(\ledr|data_out[15]~q ),
	.data_out_16(\ledr|data_out[16]~q ),
	.data_out_17(\ledr|data_out[17]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios2_qsys_0|cpu|d_writedata[17]~q ,\nios2_qsys_0|cpu|d_writedata[16]~q ,\nios2_qsys_0|cpu|d_writedata[15]~q ,\nios2_qsys_0|cpu|d_writedata[14]~q ,\nios2_qsys_0|cpu|d_writedata[13]~q ,
\nios2_qsys_0|cpu|d_writedata[12]~q ,\nios2_qsys_0|cpu|d_writedata[11]~q ,\nios2_qsys_0|cpu|d_writedata[10]~q ,\nios2_qsys_0|cpu|d_writedata[9]~q ,\nios2_qsys_0|cpu|d_writedata[8]~q ,\nios2_qsys_0|cpu|d_writedata[7]~q ,\nios2_qsys_0|cpu|d_writedata[6]~q ,
\nios2_qsys_0|cpu|d_writedata[5]~q ,\nios2_qsys_0|cpu|d_writedata[4]~q ,\nios2_qsys_0|cpu|d_writedata[3]~q ,\nios2_qsys_0|cpu|d_writedata[2]~q ,\nios2_qsys_0|cpu|d_writedata[1]~q ,\nios2_qsys_0|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.always0(\ledg|always0~1_combout ),
	.Equal2(\mm_interconnect_0|router|Equal2~1_combout ),
	.mem_used_1(\mm_interconnect_0|ledr_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always01(\ledr|always0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|ledr_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|ledr_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\ledr|readdata[0]~combout ),
	.readdata_1(\ledr|readdata[1]~combout ),
	.readdata_2(\ledr|readdata[2]~combout ),
	.readdata_3(\ledr|readdata[3]~combout ),
	.readdata_4(\ledr|readdata[4]~combout ),
	.readdata_5(\ledr|readdata[5]~combout ),
	.readdata_6(\ledr|readdata[6]~combout ),
	.readdata_7(\ledr|readdata[7]~combout ),
	.readdata_8(\ledr|readdata[8]~combout ),
	.readdata_9(\ledr|readdata[9]~combout ),
	.readdata_10(\ledr|readdata[10]~combout ),
	.readdata_11(\ledr|readdata[11]~combout ),
	.readdata_12(\ledr|readdata[12]~combout ),
	.readdata_13(\ledr|readdata[13]~combout ),
	.readdata_14(\ledr|readdata[14]~combout ),
	.readdata_15(\ledr|readdata[15]~combout ),
	.readdata_16(\ledr|readdata[16]~combout ),
	.readdata_17(\ledr|readdata[17]~combout ),
	.clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_LEDG ledg(
	.W_alu_result_7(\nios2_qsys_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_5(\nios2_qsys_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_2(\nios2_qsys_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_qsys_0|cpu|W_alu_result[3]~q ),
	.data_out_0(\ledg|data_out[0]~q ),
	.data_out_1(\ledg|data_out[1]~q ),
	.data_out_2(\ledg|data_out[2]~q ),
	.data_out_3(\ledg|data_out[3]~q ),
	.data_out_4(\ledg|data_out[4]~q ),
	.data_out_5(\ledg|data_out[5]~q ),
	.data_out_6(\ledg|data_out[6]~q ),
	.data_out_7(\ledg|data_out[7]~q ),
	.d_write(\nios2_qsys_0|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_qsys_0_data_master_translator|write_accepted~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios2_qsys_0|cpu|d_writedata[7]~q ,\nios2_qsys_0|cpu|d_writedata[6]~q ,\nios2_qsys_0|cpu|d_writedata[5]~q ,\nios2_qsys_0|cpu|d_writedata[4]~q ,\nios2_qsys_0|cpu|d_writedata[3]~q ,
\nios2_qsys_0|cpu|d_writedata[2]~q ,\nios2_qsys_0|cpu|d_writedata[1]~q ,\nios2_qsys_0|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.Equal0(\mm_interconnect_0|router|Equal0~2_combout ),
	.mem_used_1(\mm_interconnect_0|ledg_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\ledg|always0~0_combout ),
	.always01(\ledg|always0~1_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|ledg_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|ledg_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\ledg|readdata[0]~combout ),
	.readdata_1(\ledg|readdata[1]~combout ),
	.readdata_2(\ledg|readdata[2]~combout ),
	.readdata_3(\ledg|readdata[3]~combout ),
	.readdata_4(\ledg|readdata[4]~combout ),
	.readdata_5(\ledg|readdata[5]~combout ),
	.readdata_6(\ledg|readdata[6]~combout ),
	.readdata_7(\ledg|readdata[7]~combout ),
	.clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_nios2_qsys_0 nios2_qsys_0(
	.sr_0(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[0]~q ),
	.W_alu_result_28(\nios2_qsys_0|cpu|W_alu_result[28]~q ),
	.W_alu_result_27(\nios2_qsys_0|cpu|W_alu_result[27]~q ),
	.W_alu_result_26(\nios2_qsys_0|cpu|W_alu_result[26]~q ),
	.W_alu_result_25(\nios2_qsys_0|cpu|W_alu_result[25]~q ),
	.W_alu_result_24(\nios2_qsys_0|cpu|W_alu_result[24]~q ),
	.W_alu_result_23(\nios2_qsys_0|cpu|W_alu_result[23]~q ),
	.W_alu_result_22(\nios2_qsys_0|cpu|W_alu_result[22]~q ),
	.W_alu_result_21(\nios2_qsys_0|cpu|W_alu_result[21]~q ),
	.W_alu_result_20(\nios2_qsys_0|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\nios2_qsys_0|cpu|W_alu_result[19]~q ),
	.W_alu_result_18(\nios2_qsys_0|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\nios2_qsys_0|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\nios2_qsys_0|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\nios2_qsys_0|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios2_qsys_0|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios2_qsys_0|cpu|W_alu_result[13]~q ),
	.W_alu_result_6(\nios2_qsys_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_7(\nios2_qsys_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_5(\nios2_qsys_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_4(\nios2_qsys_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_12(\nios2_qsys_0|cpu|W_alu_result[12]~q ),
	.W_alu_result_10(\nios2_qsys_0|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios2_qsys_0|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios2_qsys_0|cpu|W_alu_result[8]~q ),
	.W_alu_result_11(\nios2_qsys_0|cpu|W_alu_result[11]~q ),
	.W_alu_result_2(\nios2_qsys_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_qsys_0|cpu|W_alu_result[3]~q ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.readdata_0(\audio_config|readdata[0]~q ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.readdata_1(\audio_config|readdata[1]~q ),
	.readdata_2(\audio_config|readdata[2]~q ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.readdata_17(\audio_config|readdata[17]~q ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.readdata_8(\audio_config|readdata[8]~q ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.readdata_01(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[0]~q ),
	.readdata_11(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[1]~q ),
	.readdata_21(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[3]~q ),
	.d_writedata_31(\nios2_qsys_0|cpu|d_writedata[31]~q ),
	.d_writedata_30(\nios2_qsys_0|cpu|d_writedata[30]~q ),
	.d_writedata_29(\nios2_qsys_0|cpu|d_writedata[29]~q ),
	.d_writedata_28(\nios2_qsys_0|cpu|d_writedata[28]~q ),
	.d_writedata_27(\nios2_qsys_0|cpu|d_writedata[27]~q ),
	.d_writedata_26(\nios2_qsys_0|cpu|d_writedata[26]~q ),
	.d_writedata_25(\nios2_qsys_0|cpu|d_writedata[25]~q ),
	.d_writedata_24(\nios2_qsys_0|cpu|d_writedata[24]~q ),
	.ir_out_0(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|ir_out[1]~q ),
	.d_read(\nios2_qsys_0|cpu|d_read~q ),
	.d_write(\nios2_qsys_0|cpu|d_write~q ),
	.F_pc_26(\nios2_qsys_0|cpu|F_pc[26]~q ),
	.F_pc_25(\nios2_qsys_0|cpu|F_pc[25]~q ),
	.F_pc_24(\nios2_qsys_0|cpu|F_pc[24]~q ),
	.F_pc_23(\nios2_qsys_0|cpu|F_pc[23]~q ),
	.F_pc_22(\nios2_qsys_0|cpu|F_pc[22]~q ),
	.F_pc_21(\nios2_qsys_0|cpu|F_pc[21]~q ),
	.F_pc_20(\nios2_qsys_0|cpu|F_pc[20]~q ),
	.F_pc_19(\nios2_qsys_0|cpu|F_pc[19]~q ),
	.F_pc_18(\nios2_qsys_0|cpu|F_pc[18]~q ),
	.F_pc_17(\nios2_qsys_0|cpu|F_pc[17]~q ),
	.F_pc_16(\nios2_qsys_0|cpu|F_pc[16]~q ),
	.F_pc_15(\nios2_qsys_0|cpu|F_pc[15]~q ),
	.F_pc_14(\nios2_qsys_0|cpu|F_pc[14]~q ),
	.F_pc_13(\nios2_qsys_0|cpu|F_pc[13]~q ),
	.F_pc_12(\nios2_qsys_0|cpu|F_pc[12]~q ),
	.F_pc_11(\nios2_qsys_0|cpu|F_pc[11]~q ),
	.F_pc_10(\nios2_qsys_0|cpu|F_pc[10]~q ),
	.F_pc_8(\nios2_qsys_0|cpu|F_pc[8]~q ),
	.F_pc_7(\nios2_qsys_0|cpu|F_pc[7]~q ),
	.F_pc_6(\nios2_qsys_0|cpu|F_pc[6]~q ),
	.F_pc_5(\nios2_qsys_0|cpu|F_pc[5]~q ),
	.F_pc_3(\nios2_qsys_0|cpu|F_pc[3]~q ),
	.i_read(\nios2_qsys_0|cpu|i_read~q ),
	.F_pc_2(\nios2_qsys_0|cpu|F_pc[2]~q ),
	.F_pc_4(\nios2_qsys_0|cpu|F_pc[4]~q ),
	.F_pc_9(\nios2_qsys_0|cpu|F_pc[9]~q ),
	.d_writedata_0(\nios2_qsys_0|cpu|d_writedata[0]~q ),
	.d_byteenable_0(\nios2_qsys_0|cpu|d_byteenable[0]~q ),
	.F_pc_0(\nios2_qsys_0|cpu|F_pc[0]~q ),
	.F_pc_1(\nios2_qsys_0|cpu|F_pc[1]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_writedata_1(\nios2_qsys_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_qsys_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_qsys_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_qsys_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_qsys_0|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2_qsys_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_qsys_0|cpu|d_writedata[7]~q ),
	.d_writedata_8(\nios2_qsys_0|cpu|d_writedata[8]~q ),
	.d_writedata_9(\nios2_qsys_0|cpu|d_writedata[9]~q ),
	.d_writedata_10(\nios2_qsys_0|cpu|d_writedata[10]~q ),
	.d_writedata_11(\nios2_qsys_0|cpu|d_writedata[11]~q ),
	.d_writedata_12(\nios2_qsys_0|cpu|d_writedata[12]~q ),
	.d_writedata_13(\nios2_qsys_0|cpu|d_writedata[13]~q ),
	.d_writedata_14(\nios2_qsys_0|cpu|d_writedata[14]~q ),
	.d_writedata_15(\nios2_qsys_0|cpu|d_writedata[15]~q ),
	.d_writedata_16(\nios2_qsys_0|cpu|d_writedata[16]~q ),
	.d_writedata_17(\nios2_qsys_0|cpu|d_writedata[17]~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|audio_config_avalon_av_config_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.out_valid(\mm_interconnect_0|crosser_004|clock_xer|out_valid~combout ),
	.out_data_toggle_flopped(\mm_interconnect_0|crosser_006|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\mm_interconnect_0|crosser_006|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid1(\mm_interconnect_0|crosser_006|clock_xer|out_valid~combout ),
	.read_latency_shift_reg_02(\mm_interconnect_0|ledg_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\mm_interconnect_0|ledr_s1_translator|read_latency_shift_reg[0]~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ),
	.read_latency_shift_reg_04(\mm_interconnect_0|sdram_pll_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_01(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_01(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid3(\mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ),
	.src0_valid4(\mm_interconnect_0|rsp_demux_009|src0_valid~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.mem_67_0(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_01(\mm_interconnect_0|sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_02(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_03(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_04(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_05(\mm_interconnect_0|ledr_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_06(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][67]~q ),
	.out_data_buffer_67(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_671(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[67]~q ),
	.mem_67_07(\mm_interconnect_0|ledg_s1_agent_rsp_fifo|mem[0][67]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.debug_mem_slave_waitrequest(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_translator|av_waitrequest~2_combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_004|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_009|src1_valid~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.out_valid2(\mm_interconnect_0|crosser_005|clock_xer|out_valid~combout ),
	.out_valid3(\mm_interconnect_0|crosser_007|clock_xer|out_valid~combout ),
	.av_readdatavalid(\mm_interconnect_0|nios2_qsys_0_instruction_master_agent|av_readdatavalid~4_combout ),
	.WideOr11(\mm_interconnect_0|cmd_mux_004|WideOr1~combout ),
	.local_read(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent|local_read~0_combout ),
	.hbreak_enabled(\nios2_qsys_0|cpu|hbreak_enabled~q ),
	.av_readdata_pre_30(\mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~2_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\mm_interconnect_0|sdram_pll_pll_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_01(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[0]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|sdram_pll_pll_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_11(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_21(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.readdata_31(\audio_config|readdata[3]~q ),
	.out_data_buffer_3(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_31(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[3]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.readdata_4(\audio_config|readdata[4]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_41(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[4]~q ),
	.d_byteenable_2(\nios2_qsys_0|cpu|d_byteenable[2]~q ),
	.mem(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem~4_combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_004|src_data[46]~combout ),
	.av_readdata_pre_111(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_111(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_112(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[11]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.out_data_buffer_13(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_131(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[13]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~3_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.out_data_buffer_16(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_161(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[16]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_121(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[12]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_5(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_51(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_14(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_141(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.out_data_buffer_15(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_151(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[15]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.out_data_buffer_211(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_212(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_18(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.out_data_buffer_181(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.out_data_buffer_17(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_171(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[17]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.out_data_buffer_311(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_312(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_30(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.out_data_buffer_301(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.out_data_buffer_29(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_291(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_28(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.out_data_buffer_281(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.out_data_buffer_27(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_271(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_26(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.out_data_buffer_261(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.out_data_buffer_25(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_251(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[10]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_101(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_24(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.out_data_buffer_241(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_9(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_91(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[9]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.out_data_buffer_23(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_231(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_8(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_81(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_22(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[22]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.out_data_buffer_221(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[22]~q ),
	.readdata_7(\audio_config|readdata[7]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[7]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_71(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[7]~q ),
	.readdata_6(\audio_config|readdata[6]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_61(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[6]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.out_data_buffer_20(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_201(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[20]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.out_data_buffer_19(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_191(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[19]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~9_combout ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.dreg_1(\irq_synchronizer|sync|sync[0].u|dreg[1]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.readdata_41(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[4]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~11_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[1]~14_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~16_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~19_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~21_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[3]~24_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~26_combout ),
	.src_data_41(\mm_interconnect_0|rsp_mux|src_data[4]~29_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~32_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~35_combout ),
	.src_data_61(\mm_interconnect_0|rsp_mux|src_data[6]~38_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~41_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~combout ),
	.d_byteenable_1(\nios2_qsys_0|cpu|d_byteenable[1]~q ),
	.d_byteenable_3(\nios2_qsys_0|cpu|d_byteenable[3]~q ),
	.readdata_111(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[11]~q ),
	.readdata_13(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[13]~q ),
	.readdata_16(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[16]~q ),
	.readdata_12(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[12]~q ),
	.readdata_5(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[5]~q ),
	.readdata_14(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[14]~q ),
	.readdata_15(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[15]~q ),
	.out_data_buffer_282(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_283(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[28]~q ),
	.readdata_211(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[21]~q ),
	.d_writedata_21(\nios2_qsys_0|cpu|d_writedata[21]~q ),
	.d_writedata_18(\nios2_qsys_0|cpu|d_writedata[18]~q ),
	.readdata_18(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[18]~q ),
	.out_data_buffer_272(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_273(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[27]~q ),
	.readdata_171(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[17]~q ),
	.readdata_311(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[31]~q ),
	.out_data_buffer_262(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[26]~q ),
	.out_data_buffer_263(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[26]~q ),
	.readdata_30(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[30]~q ),
	.out_data_buffer_252(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_253(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[25]~q ),
	.readdata_29(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[29]~q ),
	.out_data_buffer_242(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[24]~q ),
	.out_data_buffer_243(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[24]~q ),
	.readdata_28(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[28]~q ),
	.src_data_23(\mm_interconnect_0|rsp_mux|src_data[23]~73_combout ),
	.readdata_27(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[27]~q ),
	.src_data_22(\mm_interconnect_0|rsp_mux|src_data[22]~combout ),
	.readdata_26(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[26]~q ),
	.src_data_211(\mm_interconnect_0|rsp_mux|src_data[21]~combout ),
	.readdata_25(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[25]~q ),
	.src_data_20(\mm_interconnect_0|rsp_mux|src_data[20]~combout ),
	.readdata_10(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[10]~q ),
	.readdata_24(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[24]~q ),
	.src_data_19(\mm_interconnect_0|rsp_mux|src_data[19]~combout ),
	.readdata_9(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[9]~q ),
	.d_writedata_23(\nios2_qsys_0|cpu|d_writedata[23]~q ),
	.readdata_23(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[23]~q ),
	.src_data_18(\mm_interconnect_0|rsp_mux|src_data[18]~combout ),
	.readdata_81(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_22(\nios2_qsys_0|cpu|d_writedata[22]~q ),
	.readdata_22(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[22]~q ),
	.readdata_71(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[7]~q ),
	.readdata_61(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[6]~q ),
	.readdata_20(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[20]~q ),
	.d_writedata_20(\nios2_qsys_0|cpu|d_writedata[20]~q ),
	.readdata_19(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[19]~q ),
	.d_writedata_19(\nios2_qsys_0|cpu|d_writedata[19]~q ),
	.src_payload7(\mm_interconnect_0|cmd_mux_004|src_payload~0_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_004|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_004|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_004|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_004|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_004|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_004|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_004|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_004|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_004|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_004|src_data[32]~combout ),
	.out_data_buffer_313(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_314(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_302(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_303(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_292(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_293(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[29]~q ),
	.src_payload9(\mm_interconnect_0|cmd_mux_004|src_payload~2_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_004|src_payload~3_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_004|src_payload~4_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_004|src_payload~5_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_004|src_payload~6_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_004|src_data[33]~combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_004|src_payload~7_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_004|src_payload~8_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_004|src_data[34]~combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_004|src_payload~9_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_004|src_payload~10_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_004|src_payload~11_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_004|src_payload~12_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_004|src_payload~13_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_004|src_payload~14_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_004|src_payload~15_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_004|src_payload~16_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_004|src_data[35]~combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_004|src_payload~17_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_004|src_payload~18_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_004|src_payload~19_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_004|src_payload~20_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_004|src_payload~21_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_004|src_payload~22_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_004|src_payload~23_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_004|src_payload~24_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_004|src_payload~25_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_004|src_payload~26_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_004|src_payload~27_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_004|src_payload~28_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_004|src_payload~29_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_004|src_payload~30_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_004|src_payload~31_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_004|src_payload~32_combout ),
	.av_ld_getting_data(\nios2_qsys_0|cpu|av_ld_getting_data~9_combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux|src_data[5]~84_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux|src_data[7]~85_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_jtag_uart_0 jtag_uart_0(
	.W_alu_result_2(\nios2_qsys_0|cpu|W_alu_result[2]~q ),
	.tdo(\jtag_uart_0|final_project_soc_jtag_uart_0_alt_jtag_atlantic|tdo~q ),
	.d_read(\nios2_qsys_0|cpu|d_read~q ),
	.d_write(\nios2_qsys_0|cpu|d_write~q ),
	.read_accepted(\mm_interconnect_0|nios2_qsys_0_data_master_translator|read_accepted~q ),
	.write_accepted(\mm_interconnect_0|nios2_qsys_0_data_master_translator|write_accepted~q ),
	.cp_valid(\mm_interconnect_0|nios2_qsys_0_data_master_agent|cp_valid~combout ),
	.uav_write(\mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_write~0_combout ),
	.d_writedata_0(\nios2_qsys_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_writedata_1(\nios2_qsys_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_qsys_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_qsys_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_qsys_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_qsys_0|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2_qsys_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_qsys_0|cpu|d_writedata[7]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~1_combout ),
	.d_writedata_10(\nios2_qsys_0|cpu|d_writedata[10]~q ),
	.uav_read(\mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_read~0_combout ),
	.rst1(\jtag_uart_0|final_project_soc_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.Equal21(\mm_interconnect_0|router|Equal2~4_combout ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.b_full(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.read_01(\jtag_uart_0|read_0~q ),
	.av_readdata_0(\jtag_uart_0|av_readdata[0]~1_combout ),
	.counter_reg_bit_3(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.b_full1(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.b_non_empty(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_31(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_21(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_01(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_11(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_41(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_51(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.av_readdata_1(\jtag_uart_0|av_readdata[1]~2_combout ),
	.av_readdata_2(\jtag_uart_0|av_readdata[2]~3_combout ),
	.av_readdata_3(\jtag_uart_0|av_readdata[3]~4_combout ),
	.av_readdata_4(\jtag_uart_0|av_readdata[4]~5_combout ),
	.av_readdata_5(\jtag_uart_0|av_readdata[5]~6_combout ),
	.av_readdata_6(\jtag_uart_0|av_readdata[6]~7_combout ),
	.av_readdata_7(\jtag_uart_0|av_readdata[7]~8_combout ),
	.ac1(\jtag_uart_0|ac~q ),
	.woverflow1(\jtag_uart_0|woverflow~q ),
	.rvalid1(\jtag_uart_0|rvalid~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_audio_pll_0 audio_pll_0(
	.locked(\audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|locked ),
	.clk_0(\audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|clk[0] ),
	.clk_clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_audio_config audio_config(
	.readdata_0(\audio_config|readdata[0]~q ),
	.readdata_1(\audio_config|readdata[1]~q ),
	.readdata_2(\audio_config|readdata[2]~q ),
	.readdata_16(\audio_config|readdata[16]~q ),
	.readdata_17(\audio_config|readdata[17]~q ),
	.readdata_8(\audio_config|readdata[8]~q ),
	.I2C_SCLK(\audio_config|Serial_Bus_Controller|serial_clk~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_001|saved_grant[1]~q ),
	.d_write(\nios2_qsys_0|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_qsys_0_data_master_translator|write_accepted~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_001|src_valid~1_combout ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.uav_write(\mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_write~0_combout ),
	.mem_used_1(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem_used[1]~q ),
	.internal_reset(\audio_config|internal_reset~2_combout ),
	.d_writedata_0(\nios2_qsys_0|cpu|d_writedata[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_writedata_1(\nios2_qsys_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_qsys_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_qsys_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_qsys_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_qsys_0|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2_qsys_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_qsys_0|cpu|d_writedata[7]~q ),
	.d_writedata_8(\nios2_qsys_0|cpu|d_writedata[8]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_001|WideOr1~combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_001|src_data[68]~combout ),
	.waitrequest1(\audio_config|waitrequest~1_combout ),
	.Equal2(\audio_config|Equal2~0_combout ),
	.s_serial_transferSTATE_1_PRE_WRITE(\audio_config|s_serial_transfer.STATE_1_PRE_WRITE~q ),
	.waitrequest2(\audio_config|waitrequest~combout ),
	.I2C_SDAT(\audio_config|Serial_Bus_Controller|serial_data~1_combout ),
	.serial_data(\audio_config|Serial_Bus_Controller|serial_data~2_combout ),
	.m0_read(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent|m0_read~combout ),
	.readdata_3(\audio_config|readdata[3]~q ),
	.readdata_4(\audio_config|readdata[4]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.d_byteenable_2(\nios2_qsys_0|cpu|d_byteenable[2]~q ),
	.src_payload1(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.readdata_5(\audio_config|readdata[5]~q ),
	.readdata_7(\audio_config|readdata[7]~q ),
	.readdata_6(\audio_config|readdata[6]~q ),
	.d_byteenable_1(\nios2_qsys_0|cpu|d_byteenable[1]~q ),
	.audio_config_wire_SDAT(\audio_config_wire_SDAT~input_o ),
	.clk_clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_mm_interconnect_0 mm_interconnect_0(
	.wire_pll7_clk_0(\sdram_pll|sd1|wire_pll7_clk[0] ),
	.W_alu_result_28(\nios2_qsys_0|cpu|W_alu_result[28]~q ),
	.W_alu_result_27(\nios2_qsys_0|cpu|W_alu_result[27]~q ),
	.W_alu_result_26(\nios2_qsys_0|cpu|W_alu_result[26]~q ),
	.W_alu_result_25(\nios2_qsys_0|cpu|W_alu_result[25]~q ),
	.W_alu_result_24(\nios2_qsys_0|cpu|W_alu_result[24]~q ),
	.W_alu_result_23(\nios2_qsys_0|cpu|W_alu_result[23]~q ),
	.W_alu_result_22(\nios2_qsys_0|cpu|W_alu_result[22]~q ),
	.W_alu_result_21(\nios2_qsys_0|cpu|W_alu_result[21]~q ),
	.W_alu_result_20(\nios2_qsys_0|cpu|W_alu_result[20]~q ),
	.W_alu_result_19(\nios2_qsys_0|cpu|W_alu_result[19]~q ),
	.W_alu_result_18(\nios2_qsys_0|cpu|W_alu_result[18]~q ),
	.W_alu_result_17(\nios2_qsys_0|cpu|W_alu_result[17]~q ),
	.W_alu_result_16(\nios2_qsys_0|cpu|W_alu_result[16]~q ),
	.W_alu_result_15(\nios2_qsys_0|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios2_qsys_0|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios2_qsys_0|cpu|W_alu_result[13]~q ),
	.W_alu_result_6(\nios2_qsys_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_7(\nios2_qsys_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_5(\nios2_qsys_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_4(\nios2_qsys_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_12(\nios2_qsys_0|cpu|W_alu_result[12]~q ),
	.W_alu_result_10(\nios2_qsys_0|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios2_qsys_0|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios2_qsys_0|cpu|W_alu_result[8]~q ),
	.W_alu_result_11(\nios2_qsys_0|cpu|W_alu_result[11]~q ),
	.W_alu_result_2(\nios2_qsys_0|cpu|W_alu_result[2]~q ),
	.W_alu_result_3(\nios2_qsys_0|cpu|W_alu_result[3]~q ),
	.clk_0(\audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|clk[0] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.readdata_0(\audio_config|readdata[0]~q ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.readdata_1(\audio_config|readdata[1]~q ),
	.readdata_2(\audio_config|readdata[2]~q ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.readdata_16(\audio_config|readdata[16]~q ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.readdata_17(\audio_config|readdata[17]~q ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.readdata_8(\audio_config|readdata[8]~q ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.readdata_01(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[0]~q ),
	.readdata_11(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[1]~q ),
	.readdata_21(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[3]~q ),
	.d_writedata_31(\nios2_qsys_0|cpu|d_writedata[31]~q ),
	.d_writedata_30(\nios2_qsys_0|cpu|d_writedata[30]~q ),
	.d_writedata_29(\nios2_qsys_0|cpu|d_writedata[29]~q ),
	.d_writedata_28(\nios2_qsys_0|cpu|d_writedata[28]~q ),
	.d_writedata_27(\nios2_qsys_0|cpu|d_writedata[27]~q ),
	.d_writedata_26(\nios2_qsys_0|cpu|d_writedata[26]~q ),
	.d_writedata_25(\nios2_qsys_0|cpu|d_writedata[25]~q ),
	.d_writedata_24(\nios2_qsys_0|cpu|d_writedata[24]~q ),
	.readdata_02(\audio|readdata[0]~q ),
	.readdata_12(\audio|readdata[1]~q ),
	.readdata_22(\audio|readdata[2]~q ),
	.readdata_31(\audio|readdata[3]~q ),
	.readdata_4(\audio|readdata[4]~q ),
	.readdata_111(\audio|readdata[11]~q ),
	.readdata_13(\audio|readdata[13]~q ),
	.readdata_161(\audio|readdata[16]~q ),
	.readdata_121(\audio|readdata[12]~q ),
	.readdata_5(\audio|readdata[5]~q ),
	.readdata_14(\audio|readdata[14]~q ),
	.readdata_15(\audio|readdata[15]~q ),
	.readdata_211(\audio|readdata[21]~q ),
	.readdata_18(\audio|readdata[18]~q ),
	.readdata_171(\audio|readdata[17]~q ),
	.readdata_311(\audio|readdata[31]~q ),
	.readdata_30(\audio|readdata[30]~q ),
	.readdata_29(\audio|readdata[29]~q ),
	.readdata_28(\audio|readdata[28]~q ),
	.readdata_27(\audio|readdata[27]~q ),
	.readdata_26(\audio|readdata[26]~q ),
	.readdata_25(\audio|readdata[25]~q ),
	.readdata_10(\audio|readdata[10]~q ),
	.readdata_24(\audio|readdata[24]~q ),
	.readdata_9(\audio|readdata[9]~q ),
	.readdata_23(\audio|readdata[23]~q ),
	.readdata_81(\audio|readdata[8]~q ),
	.readdata_221(\audio|readdata[22]~q ),
	.readdata_7(\audio|readdata[7]~q ),
	.readdata_6(\audio|readdata[6]~q ),
	.readdata_20(\audio|readdata[20]~q ),
	.readdata_19(\audio|readdata[19]~q ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_001|saved_grant[1]~q ),
	.d_read(\nios2_qsys_0|cpu|d_read~q ),
	.d_write(\nios2_qsys_0|cpu|d_write~q ),
	.read_accepted(\mm_interconnect_0|nios2_qsys_0_data_master_translator|read_accepted~q ),
	.write_accepted(\mm_interconnect_0|nios2_qsys_0_data_master_translator|write_accepted~q ),
	.cp_valid(\mm_interconnect_0|nios2_qsys_0_data_master_agent|cp_valid~combout ),
	.src_valid(\mm_interconnect_0|cmd_mux_001|src_valid~1_combout ),
	.F_pc_26(\nios2_qsys_0|cpu|F_pc[26]~q ),
	.F_pc_25(\nios2_qsys_0|cpu|F_pc[25]~q ),
	.F_pc_24(\nios2_qsys_0|cpu|F_pc[24]~q ),
	.F_pc_23(\nios2_qsys_0|cpu|F_pc[23]~q ),
	.F_pc_22(\nios2_qsys_0|cpu|F_pc[22]~q ),
	.F_pc_21(\nios2_qsys_0|cpu|F_pc[21]~q ),
	.F_pc_20(\nios2_qsys_0|cpu|F_pc[20]~q ),
	.F_pc_19(\nios2_qsys_0|cpu|F_pc[19]~q ),
	.F_pc_18(\nios2_qsys_0|cpu|F_pc[18]~q ),
	.F_pc_17(\nios2_qsys_0|cpu|F_pc[17]~q ),
	.F_pc_16(\nios2_qsys_0|cpu|F_pc[16]~q ),
	.F_pc_15(\nios2_qsys_0|cpu|F_pc[15]~q ),
	.F_pc_14(\nios2_qsys_0|cpu|F_pc[14]~q ),
	.F_pc_13(\nios2_qsys_0|cpu|F_pc[13]~q ),
	.F_pc_12(\nios2_qsys_0|cpu|F_pc[12]~q ),
	.F_pc_11(\nios2_qsys_0|cpu|F_pc[11]~q ),
	.F_pc_10(\nios2_qsys_0|cpu|F_pc[10]~q ),
	.F_pc_8(\nios2_qsys_0|cpu|F_pc[8]~q ),
	.F_pc_7(\nios2_qsys_0|cpu|F_pc[7]~q ),
	.F_pc_6(\nios2_qsys_0|cpu|F_pc[6]~q ),
	.F_pc_5(\nios2_qsys_0|cpu|F_pc[5]~q ),
	.F_pc_3(\nios2_qsys_0|cpu|F_pc[3]~q ),
	.i_read(\nios2_qsys_0|cpu|i_read~q ),
	.F_pc_2(\nios2_qsys_0|cpu|F_pc[2]~q ),
	.F_pc_4(\nios2_qsys_0|cpu|F_pc[4]~q ),
	.F_pc_9(\nios2_qsys_0|cpu|F_pc[9]~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.uav_write(\mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_write~0_combout ),
	.mem_used_1(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem_used[1]~q ),
	.internal_reset(\audio_config|internal_reset~2_combout ),
	.d_writedata_0(\nios2_qsys_0|cpu|d_writedata[0]~q ),
	.d_byteenable_0(\nios2_qsys_0|cpu|d_byteenable[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.F_pc_0(\nios2_qsys_0|cpu|F_pc[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.F_pc_1(\nios2_qsys_0|cpu|F_pc[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.Equal0(\mm_interconnect_0|router|Equal0~2_combout ),
	.mem_used_11(\mm_interconnect_0|ledg_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\ledg|always0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|ledg_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|ledg_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_1(\nios2_qsys_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_qsys_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_qsys_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_qsys_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_qsys_0|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios2_qsys_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_qsys_0|cpu|d_writedata[7]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~1_combout ),
	.mem_used_12(\mm_interconnect_0|ledr_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always01(\ledr|always0~0_combout ),
	.wait_latency_counter_11(\mm_interconnect_0|ledr_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|ledr_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_8(\nios2_qsys_0|cpu|d_writedata[8]~q ),
	.d_writedata_9(\nios2_qsys_0|cpu|d_writedata[9]~q ),
	.d_writedata_10(\nios2_qsys_0|cpu|d_writedata[10]~q ),
	.d_writedata_11(\nios2_qsys_0|cpu|d_writedata[11]~q ),
	.d_writedata_12(\nios2_qsys_0|cpu|d_writedata[12]~q ),
	.d_writedata_13(\nios2_qsys_0|cpu|d_writedata[13]~q ),
	.d_writedata_14(\nios2_qsys_0|cpu|d_writedata[14]~q ),
	.d_writedata_15(\nios2_qsys_0|cpu|d_writedata[15]~q ),
	.d_writedata_16(\nios2_qsys_0|cpu|d_writedata[16]~q ),
	.d_writedata_17(\nios2_qsys_0|cpu|d_writedata[17]~q ),
	.entries_1(\sdram|the_final_project_soc_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_final_project_soc_sdram_input_efifo_module|entries[0]~q ),
	.altera_reset_synchronizer_int_chain_out1(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_001|WideOr1~combout ),
	.uav_read(\mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_read~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_001|src_data[68]~combout ),
	.waitrequest(\audio_config|waitrequest~1_combout ),
	.Equal21(\audio_config|Equal2~0_combout ),
	.s_serial_transferSTATE_1_PRE_WRITE(\audio_config|s_serial_transfer.STATE_1_PRE_WRITE~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|audio_config_avalon_av_config_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.out_valid(\mm_interconnect_0|crosser_004|clock_xer|out_valid~combout ),
	.out_data_toggle_flopped(\mm_interconnect_0|crosser_006|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\mm_interconnect_0|crosser_006|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid1(\mm_interconnect_0|crosser_006|clock_xer|out_valid~combout ),
	.read_latency_shift_reg_02(\mm_interconnect_0|ledg_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\mm_interconnect_0|ledr_s1_translator|read_latency_shift_reg[0]~q ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_003|src0_valid~0_combout ),
	.src0_valid2(\mm_interconnect_0|rsp_demux_004|src0_valid~0_combout ),
	.read_latency_shift_reg_04(\mm_interconnect_0|sdram_pll_pll_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_01(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_01(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid3(\mm_interconnect_0|rsp_demux_005|src0_valid~0_combout ),
	.src0_valid4(\mm_interconnect_0|rsp_demux_009|src0_valid~0_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.mem_67_0(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_01(\mm_interconnect_0|sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_02(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_03(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_04(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_05(\mm_interconnect_0|ledr_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_67_06(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][67]~q ),
	.out_data_buffer_67(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_671(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[67]~q ),
	.mem_67_07(\mm_interconnect_0|ledg_s1_agent_rsp_fifo|mem[0][67]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.rst1(\jtag_uart_0|final_project_soc_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.Equal22(\mm_interconnect_0|router|Equal2~4_combout ),
	.av_waitrequest(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_13(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.waitrequest1(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_14(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.mem_used_15(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_009|saved_grant[0]~q ),
	.mem_used_16(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.waitrequest2(\audio_config|waitrequest~combout ),
	.nios2_qsys_0_data_master_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_translator|av_waitrequest~2_combout ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_004|src1_valid~0_combout ),
	.src1_valid3(\mm_interconnect_0|rsp_demux_009|src1_valid~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.out_valid2(\mm_interconnect_0|crosser_005|clock_xer|out_valid~combout ),
	.out_valid3(\mm_interconnect_0|crosser_007|clock_xer|out_valid~combout ),
	.av_readdatavalid(\mm_interconnect_0|nios2_qsys_0_instruction_master_agent|av_readdatavalid~4_combout ),
	.saved_grant_02(\mm_interconnect_0|cmd_mux|saved_grant[0]~q ),
	.out_data_buffer_3(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[3]~q ),
	.src_data_381(\mm_interconnect_0|cmd_mux|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux|src_data[39]~combout ),
	.WideOr12(\mm_interconnect_0|cmd_mux|WideOr1~combout ),
	.mem_used_17(\mm_interconnect_0|audio_avalon_audio_slave_agent_rsp_fifo|mem_used[1]~q ),
	.last_cycle(\mm_interconnect_0|cmd_mux|last_cycle~0_combout ),
	.nonposted_write_endofpacket(\mm_interconnect_0|audio_avalon_audio_slave_agent|nonposted_write_endofpacket~0_combout ),
	.WideOr13(\mm_interconnect_0|cmd_mux_005|WideOr1~combout ),
	.src_data_382(\mm_interconnect_0|cmd_mux_005|src_data[38]~combout ),
	.mem(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem~0_combout ),
	.src_data_392(\mm_interconnect_0|cmd_mux_005|src_data[39]~combout ),
	.last_cycle1(\mm_interconnect_0|cmd_mux_006|last_cycle~0_combout ),
	.saved_grant_11(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.WideOr14(\mm_interconnect_0|cmd_mux_006|WideOr1~combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_006|src_payload~0_combout ),
	.src_data_681(\mm_interconnect_0|cmd_mux_006|src_data[68]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_006|src_data[48]~combout ),
	.src_data_62(\mm_interconnect_0|cmd_mux_006|src_data[62]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_006|src_data[49]~combout ),
	.src_data_51(\mm_interconnect_0|cmd_mux_006|src_data[51]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_006|src_data[50]~combout ),
	.src_data_53(\mm_interconnect_0|cmd_mux_006|src_data[53]~combout ),
	.src_data_52(\mm_interconnect_0|cmd_mux_006|src_data[52]~combout ),
	.src_data_55(\mm_interconnect_0|cmd_mux_006|src_data[55]~combout ),
	.src_data_54(\mm_interconnect_0|cmd_mux_006|src_data[54]~combout ),
	.src_data_57(\mm_interconnect_0|cmd_mux_006|src_data[57]~combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_006|src_data[56]~combout ),
	.src_data_59(\mm_interconnect_0|cmd_mux_006|src_data[59]~combout ),
	.src_data_58(\mm_interconnect_0|cmd_mux_006|src_data[58]~combout ),
	.src_data_61(\mm_interconnect_0|cmd_mux_006|src_data[61]~combout ),
	.src_data_60(\mm_interconnect_0|cmd_mux_006|src_data[60]~combout ),
	.src_data_383(\mm_interconnect_0|cmd_mux_006|src_data[38]~combout ),
	.src_data_393(\mm_interconnect_0|cmd_mux_006|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_006|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_006|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_006|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_006|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_006|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_006|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_006|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_006|src_data[47]~combout ),
	.out_data_buffer_32(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_321(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_33(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_331(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_34(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_341(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_35(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[35]~q ),
	.out_data_buffer_351(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[35]~q ),
	.m0_read(\mm_interconnect_0|audio_config_avalon_av_config_slave_agent|m0_read~combout ),
	.WideOr15(\mm_interconnect_0|cmd_mux_004|WideOr1~combout ),
	.local_read(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent|local_read~0_combout ),
	.mem1(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr16(\mm_interconnect_0|cmd_mux_009|WideOr1~combout ),
	.hbreak_enabled(\nios2_qsys_0|cpu|hbreak_enabled~q ),
	.av_readdata_pre_30(\mm_interconnect_0|sysid_qsys_0_control_slave_translator|av_readdata_pre[30]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~2_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\mm_interconnect_0|sdram_pll_pll_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_0(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_01(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[0]~q ),
	.av_readdata_pre_1(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_11(\mm_interconnect_0|sdram_pll_pll_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_11(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_21(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_3(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.readdata_32(\audio_config|readdata[3]~q ),
	.out_data_buffer_31(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_36(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[3]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.readdata_41(\audio_config|readdata[4]~q ),
	.out_data_buffer_4(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_41(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[4]~q ),
	.src_payload5(\mm_interconnect_0|cmd_mux|src_payload~0_combout ),
	.src_data_682(\mm_interconnect_0|cmd_mux|src_data[68]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.d_byteenable_2(\nios2_qsys_0|cpu|d_byteenable[2]~q ),
	.src_payload7(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.mem2(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem~4_combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_004|src_data[46]~combout ),
	.av_readdata_pre_111(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.out_data_buffer_111(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_112(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[11]~q ),
	.av_readdata_pre_13(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.out_data_buffer_13(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_131(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[13]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~3_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.out_data_buffer_16(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_161(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[16]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_121(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[12]~q ),
	.readdata_51(\audio_config|readdata[5]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_5(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_5(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_51(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_14(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_141(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_15(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.out_data_buffer_15(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_151(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[15]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.out_data_buffer_211(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_212(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_18(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.out_data_buffer_181(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.out_data_buffer_17(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_171(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[17]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.out_data_buffer_311(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_312(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_30(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.out_data_buffer_301(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[30]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.out_data_buffer_29(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_291(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_28(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.out_data_buffer_281(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[28]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.out_data_buffer_27(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_271(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_26(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.out_data_buffer_261(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[26]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.out_data_buffer_25(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_251(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_10(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[10]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_101(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_24(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.out_data_buffer_241(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[24]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_9(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_91(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[9]~q ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.out_data_buffer_23(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_231(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_8(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_81(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_22(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[22]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.out_data_buffer_221(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[22]~q ),
	.readdata_71(\audio_config|readdata[7]~q ),
	.out_data_buffer_7(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[7]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_71(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[7]~q ),
	.readdata_61(\audio_config|readdata[6]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_6(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_61(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[6]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.out_data_buffer_20(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_201(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[20]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|nios2_qsys_0_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.out_data_buffer_19(\mm_interconnect_0|crosser_007|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_191(\mm_interconnect_0|crosser_005|clock_xer|out_data_buffer[19]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~9_combout ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_009|src_payload~0_combout ),
	.src_data_384(\mm_interconnect_0|cmd_mux_009|src_data[38]~combout ),
	.src_data_394(\mm_interconnect_0|cmd_mux_009|src_data[39]~combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_009|src_data[32]~combout ),
	.readdata_03(\sdram_pll|readdata[0]~1_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_009|src_payload~1_combout ),
	.readdata_110(\sdram_pll|readdata[1]~2_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_009|src_payload~2_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_009|src_payload~3_combout ),
	.readdata_42(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[4]~q ),
	.src_payload15(\mm_interconnect_0|cmd_mux_009|src_payload~4_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux|src_payload~1_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~11_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[1]~14_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~16_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~19_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~21_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[3]~24_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~26_combout ),
	.src_data_410(\mm_interconnect_0|rsp_mux|src_data[4]~29_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~32_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~35_combout ),
	.src_data_63(\mm_interconnect_0|rsp_mux|src_data[6]~38_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~41_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~combout ),
	.d_byteenable_1(\nios2_qsys_0|cpu|d_byteenable[1]~q ),
	.d_byteenable_3(\nios2_qsys_0|cpu|d_byteenable[3]~q ),
	.b_full(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_payload17(\mm_interconnect_0|cmd_mux_006|src_payload~1_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_006|src_payload~2_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_006|src_payload~3_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_006|src_payload~4_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_006|src_payload~5_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_006|src_payload~6_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_006|src_payload~7_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_006|src_payload~8_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_006|src_payload~9_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_006|src_payload~10_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_006|src_payload~11_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_006|src_payload~12_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_006|src_payload~13_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_006|src_payload~14_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_006|src_payload~15_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_006|src_payload~16_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_006|src_payload~17_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_006|src_payload~18_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_006|src_payload~19_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_006|src_payload~20_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_006|src_payload~21_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_006|src_payload~22_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_006|src_payload~23_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_006|src_payload~24_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_006|src_payload~25_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_006|src_payload~26_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_006|src_payload~27_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_006|src_payload~28_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_006|src_payload~29_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_006|src_payload~30_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_006|src_payload~31_combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_006|src_payload~32_combout ),
	.readdata_112(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[11]~q ),
	.src_payload49(\mm_interconnect_0|cmd_mux_009|src_payload~5_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_009|src_data[33]~combout ),
	.readdata_131(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[13]~q ),
	.src_payload50(\mm_interconnect_0|cmd_mux_009|src_payload~6_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_009|src_payload~7_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_009|src_data[34]~combout ),
	.readdata_162(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[16]~q ),
	.src_payload52(\mm_interconnect_0|cmd_mux_009|src_payload~8_combout ),
	.readdata_122(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[12]~q ),
	.src_payload53(\mm_interconnect_0|cmd_mux_009|src_payload~9_combout ),
	.readdata_52(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[5]~q ),
	.src_payload54(\mm_interconnect_0|cmd_mux_009|src_payload~10_combout ),
	.readdata_141(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[14]~q ),
	.readdata_151(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[15]~q ),
	.src_payload55(\mm_interconnect_0|cmd_mux_009|src_payload~11_combout ),
	.out_data_buffer_282(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_283(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[28]~q ),
	.readdata_212(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[21]~q ),
	.d_writedata_21(\nios2_qsys_0|cpu|d_writedata[21]~q ),
	.src_payload56(\mm_interconnect_0|cmd_mux_009|src_payload~12_combout ),
	.d_writedata_18(\nios2_qsys_0|cpu|d_writedata[18]~q ),
	.src_payload57(\mm_interconnect_0|cmd_mux_009|src_payload~13_combout ),
	.readdata_181(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[18]~q ),
	.out_data_buffer_272(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_273(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[27]~q ),
	.readdata_172(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[17]~q ),
	.src_payload58(\mm_interconnect_0|cmd_mux_009|src_payload~14_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_009|src_payload~15_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_009|src_data[35]~combout ),
	.readdata_312(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[31]~q ),
	.out_data_buffer_262(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[26]~q ),
	.out_data_buffer_263(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[26]~q ),
	.src_payload60(\mm_interconnect_0|cmd_mux_009|src_payload~16_combout ),
	.readdata_301(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[30]~q ),
	.out_data_buffer_252(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_253(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[25]~q ),
	.src_payload61(\mm_interconnect_0|cmd_mux_009|src_payload~17_combout ),
	.readdata_291(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[29]~q ),
	.out_data_buffer_242(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[24]~q ),
	.out_data_buffer_243(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[24]~q ),
	.src_payload62(\mm_interconnect_0|cmd_mux_009|src_payload~18_combout ),
	.readdata_281(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[28]~q ),
	.src_data_23(\mm_interconnect_0|rsp_mux|src_data[23]~73_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_009|src_payload~19_combout ),
	.readdata_271(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[27]~q ),
	.src_data_22(\mm_interconnect_0|rsp_mux|src_data[22]~combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_009|src_payload~20_combout ),
	.readdata_261(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[26]~q ),
	.src_data_211(\mm_interconnect_0|rsp_mux|src_data[21]~combout ),
	.src_payload65(\mm_interconnect_0|cmd_mux_009|src_payload~21_combout ),
	.readdata_251(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[25]~q ),
	.src_data_20(\mm_interconnect_0|rsp_mux|src_data[20]~combout ),
	.src_payload66(\mm_interconnect_0|cmd_mux_009|src_payload~22_combout ),
	.readdata_101(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[10]~q ),
	.src_payload67(\mm_interconnect_0|cmd_mux_009|src_payload~23_combout ),
	.readdata_241(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[24]~q ),
	.src_data_19(\mm_interconnect_0|rsp_mux|src_data[19]~combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_009|src_payload~24_combout ),
	.readdata_91(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[9]~q ),
	.d_writedata_23(\nios2_qsys_0|cpu|d_writedata[23]~q ),
	.src_payload69(\mm_interconnect_0|cmd_mux_009|src_payload~25_combout ),
	.readdata_231(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[23]~q ),
	.src_data_18(\mm_interconnect_0|rsp_mux|src_data[18]~combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_009|src_payload~26_combout ),
	.readdata_82(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_22(\nios2_qsys_0|cpu|d_writedata[22]~q ),
	.src_payload71(\mm_interconnect_0|cmd_mux_009|src_payload~27_combout ),
	.readdata_222(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[22]~q ),
	.src_payload72(\mm_interconnect_0|cmd_mux_009|src_payload~28_combout ),
	.readdata_72(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[7]~q ),
	.src_payload73(\mm_interconnect_0|cmd_mux_009|src_payload~29_combout ),
	.readdata_62(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[6]~q ),
	.readdata_201(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[20]~q ),
	.d_writedata_20(\nios2_qsys_0|cpu|d_writedata[20]~q ),
	.src_payload74(\mm_interconnect_0|cmd_mux_009|src_payload~30_combout ),
	.readdata_191(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|readdata[19]~q ),
	.d_writedata_19(\nios2_qsys_0|cpu|d_writedata[19]~q ),
	.src_payload75(\mm_interconnect_0|cmd_mux_009|src_payload~31_combout ),
	.readdata_04(\ledr|readdata[0]~combout ),
	.read_0(\jtag_uart_0|read_0~q ),
	.av_readdata_0(\jtag_uart_0|av_readdata[0]~1_combout ),
	.readdata_05(\ledg|readdata[0]~combout ),
	.counter_reg_bit_3(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.b_full1(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.b_non_empty(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_31(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_21(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_01(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_11(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_41(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_51(\jtag_uart_0|the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.src_payload76(\mm_interconnect_0|cmd_mux|src_payload~2_combout ),
	.readdata_113(\ledr|readdata[1]~combout ),
	.av_readdata_1(\jtag_uart_0|av_readdata[1]~2_combout ),
	.readdata_114(\ledg|readdata[1]~combout ),
	.readdata_210(\ledr|readdata[2]~combout ),
	.av_readdata_2(\jtag_uart_0|av_readdata[2]~3_combout ),
	.readdata_213(\ledg|readdata[2]~combout ),
	.readdata_33(\ledr|readdata[3]~combout ),
	.av_readdata_3(\jtag_uart_0|av_readdata[3]~4_combout ),
	.readdata_34(\ledg|readdata[3]~combout ),
	.readdata_43(\ledr|readdata[4]~combout ),
	.av_readdata_4(\jtag_uart_0|av_readdata[4]~5_combout ),
	.readdata_44(\ledg|readdata[4]~combout ),
	.readdata_53(\ledr|readdata[5]~combout ),
	.av_readdata_5(\jtag_uart_0|av_readdata[5]~6_combout ),
	.readdata_54(\ledg|readdata[5]~combout ),
	.readdata_63(\ledr|readdata[6]~combout ),
	.av_readdata_6(\jtag_uart_0|av_readdata[6]~7_combout ),
	.readdata_64(\ledg|readdata[6]~combout ),
	.readdata_73(\ledr|readdata[7]~combout ),
	.av_readdata_7(\jtag_uart_0|av_readdata[7]~8_combout ),
	.readdata_74(\ledg|readdata[7]~combout ),
	.readdata_83(\ledr|readdata[8]~combout ),
	.readdata_92(\ledr|readdata[9]~combout ),
	.readdata_102(\ledr|readdata[10]~combout ),
	.ac(\jtag_uart_0|ac~q ),
	.readdata_115(\ledr|readdata[11]~combout ),
	.readdata_123(\ledr|readdata[12]~combout ),
	.readdata_132(\ledr|readdata[13]~combout ),
	.readdata_142(\ledr|readdata[14]~combout ),
	.woverflow(\jtag_uart_0|woverflow~q ),
	.readdata_152(\ledr|readdata[15]~combout ),
	.rvalid(\jtag_uart_0|rvalid~q ),
	.readdata_163(\ledr|readdata[16]~combout ),
	.readdata_173(\ledr|readdata[17]~combout ),
	.src_payload77(\mm_interconnect_0|cmd_mux_004|src_payload~0_combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_004|src_payload~1_combout ),
	.src_data_385(\mm_interconnect_0|cmd_mux_004|src_data[38]~combout ),
	.src_data_395(\mm_interconnect_0|cmd_mux_004|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_004|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_004|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_004|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_004|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_004|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_004|src_data[45]~combout ),
	.src_data_322(\mm_interconnect_0|cmd_mux_004|src_data[32]~combout ),
	.out_data_buffer_313(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_314(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_302(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_303(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_292(\mm_interconnect_0|crosser_006|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_293(\mm_interconnect_0|crosser_004|clock_xer|out_data_buffer[29]~q ),
	.src_payload79(\mm_interconnect_0|cmd_mux_004|src_payload~2_combout ),
	.src_payload80(\mm_interconnect_0|cmd_mux_004|src_payload~3_combout ),
	.src_payload81(\mm_interconnect_0|cmd_mux|src_payload~3_combout ),
	.za_valid(\sdram|za_valid~q ),
	.out_data_buffer_02(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_110(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[1]~q ),
	.src_payload82(\mm_interconnect_0|cmd_mux_004|src_payload~4_combout ),
	.out_data_buffer_210(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[2]~q ),
	.src_payload83(\mm_interconnect_0|cmd_mux_004|src_payload~5_combout ),
	.src_payload84(\mm_interconnect_0|cmd_mux|src_payload~4_combout ),
	.src_payload85(\mm_interconnect_0|cmd_mux_004|src_payload~6_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_004|src_data[33]~combout ),
	.src_payload86(\mm_interconnect_0|cmd_mux_004|src_payload~7_combout ),
	.src_payload87(\mm_interconnect_0|cmd_mux_004|src_payload~8_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_004|src_data[34]~combout ),
	.src_payload88(\mm_interconnect_0|cmd_mux_004|src_payload~9_combout ),
	.src_payload89(\mm_interconnect_0|cmd_mux_004|src_payload~10_combout ),
	.src_payload90(\mm_interconnect_0|cmd_mux_004|src_payload~11_combout ),
	.src_payload91(\mm_interconnect_0|cmd_mux_004|src_payload~12_combout ),
	.src_payload92(\mm_interconnect_0|cmd_mux_004|src_payload~13_combout ),
	.src_payload93(\mm_interconnect_0|cmd_mux_004|src_payload~14_combout ),
	.src_payload94(\mm_interconnect_0|cmd_mux_004|src_payload~15_combout ),
	.src_payload95(\mm_interconnect_0|cmd_mux_004|src_payload~16_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_004|src_data[35]~combout ),
	.src_payload96(\mm_interconnect_0|cmd_mux_004|src_payload~17_combout ),
	.src_payload97(\mm_interconnect_0|cmd_mux_004|src_payload~18_combout ),
	.src_payload98(\mm_interconnect_0|cmd_mux_004|src_payload~19_combout ),
	.src_payload99(\mm_interconnect_0|cmd_mux_004|src_payload~20_combout ),
	.src_payload100(\mm_interconnect_0|cmd_mux_004|src_payload~21_combout ),
	.src_payload101(\mm_interconnect_0|cmd_mux_004|src_payload~22_combout ),
	.src_payload102(\mm_interconnect_0|cmd_mux_004|src_payload~23_combout ),
	.src_payload103(\mm_interconnect_0|cmd_mux_004|src_payload~24_combout ),
	.src_payload104(\mm_interconnect_0|cmd_mux_004|src_payload~25_combout ),
	.src_payload105(\mm_interconnect_0|cmd_mux_004|src_payload~26_combout ),
	.src_payload106(\mm_interconnect_0|cmd_mux_004|src_payload~27_combout ),
	.src_payload107(\mm_interconnect_0|cmd_mux_004|src_payload~28_combout ),
	.src_payload108(\mm_interconnect_0|cmd_mux_004|src_payload~29_combout ),
	.src_payload109(\mm_interconnect_0|cmd_mux_004|src_payload~30_combout ),
	.src_payload110(\mm_interconnect_0|cmd_mux_004|src_payload~31_combout ),
	.src_payload111(\mm_interconnect_0|cmd_mux_004|src_payload~32_combout ),
	.za_data_0(\sdram|za_data[0]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.src_payload112(\mm_interconnect_0|cmd_mux|src_payload~5_combout ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.za_data_16(\sdram|za_data[16]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.za_data_21(\sdram|za_data[21]~q ),
	.za_data_18(\sdram|za_data[18]~q ),
	.za_data_17(\sdram|za_data[17]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.za_data_23(\sdram|za_data[23]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.za_data_22(\sdram|za_data[22]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.za_data_20(\sdram|za_data[20]~q ),
	.za_data_19(\sdram|za_data[19]~q ),
	.src_payload113(\mm_interconnect_0|cmd_mux|src_payload~6_combout ),
	.src_payload114(\mm_interconnect_0|cmd_mux|src_payload~7_combout ),
	.src_payload115(\mm_interconnect_0|cmd_mux|src_payload~8_combout ),
	.src_payload116(\mm_interconnect_0|cmd_mux|src_payload~9_combout ),
	.src_payload117(\mm_interconnect_0|cmd_mux|src_payload~10_combout ),
	.src_payload118(\mm_interconnect_0|cmd_mux|src_payload~11_combout ),
	.src_payload119(\mm_interconnect_0|cmd_mux|src_payload~12_combout ),
	.src_payload120(\mm_interconnect_0|cmd_mux|src_payload~13_combout ),
	.src_payload121(\mm_interconnect_0|cmd_mux|src_payload~14_combout ),
	.src_payload122(\mm_interconnect_0|cmd_mux|src_payload~15_combout ),
	.src_payload123(\mm_interconnect_0|cmd_mux|src_payload~16_combout ),
	.src_payload124(\mm_interconnect_0|cmd_mux|src_payload~17_combout ),
	.src_payload125(\mm_interconnect_0|cmd_mux|src_payload~18_combout ),
	.src_payload126(\mm_interconnect_0|cmd_mux|src_payload~19_combout ),
	.src_payload127(\mm_interconnect_0|cmd_mux|src_payload~20_combout ),
	.src_payload128(\mm_interconnect_0|cmd_mux|src_payload~21_combout ),
	.src_payload129(\mm_interconnect_0|cmd_mux|src_payload~22_combout ),
	.src_payload130(\mm_interconnect_0|cmd_mux|src_payload~23_combout ),
	.src_payload131(\mm_interconnect_0|cmd_mux|src_payload~24_combout ),
	.src_payload132(\mm_interconnect_0|cmd_mux|src_payload~25_combout ),
	.src_payload133(\mm_interconnect_0|cmd_mux|src_payload~26_combout ),
	.src_payload134(\mm_interconnect_0|cmd_mux|src_payload~27_combout ),
	.src_payload135(\mm_interconnect_0|cmd_mux|src_payload~28_combout ),
	.src_payload136(\mm_interconnect_0|cmd_mux|src_payload~29_combout ),
	.src_payload137(\mm_interconnect_0|cmd_mux|src_payload~30_combout ),
	.src_payload138(\mm_interconnect_0|cmd_mux|src_payload~31_combout ),
	.av_ld_getting_data(\nios2_qsys_0|cpu|av_ld_getting_data~9_combout ),
	.m0_write(\mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ),
	.src_data_510(\mm_interconnect_0|rsp_mux|src_data[5]~84_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux|src_data[7]~85_combout ),
	.clk_clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_sdram_pll sdram_pll(
	.wire_pll7_clk_0(\sdram_pll|sd1|wire_pll7_clk[0] ),
	.wire_pll7_clk_1(\sdram_pll|sd1|wire_pll7_clk[1] ),
	.locked(\sdram_pll|sd1|locked~combout ),
	.d_writedata_0(\nios2_qsys_0|cpu|d_writedata[0]~q ),
	.reset(\rst_controller|r_sync_rst~q ),
	.d_writedata_1(\nios2_qsys_0|cpu|d_writedata[1]~q ),
	.mem_used_1(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_005|WideOr1~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_005|src_data[38]~combout ),
	.mem(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem~0_combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_005|src_data[39]~combout ),
	.mem1(\mm_interconnect_0|sdram_pll_pll_slave_agent_rsp_fifo|mem~1_combout ),
	.readdata_0(\sdram_pll|readdata[0]~1_combout ),
	.readdata_1(\sdram_pll|readdata[1]~2_combout ),
	.clk_clk(\clk_clk~input_o ),
	.unused_sdram_areset_conduit_export(\unused_sdram_areset_conduit_export~input_o ));

final_project_soc_final_project_soc_sdram sdram(
	.wire_pll7_clk_0(\sdram_pll|sd1|wire_pll7_clk[0] ),
	.m_addr_0(\sdram|m_addr[0]~q ),
	.m_addr_1(\sdram|m_addr[1]~q ),
	.m_addr_2(\sdram|m_addr[2]~q ),
	.m_addr_3(\sdram|m_addr[3]~q ),
	.m_addr_4(\sdram|m_addr[4]~q ),
	.m_addr_5(\sdram|m_addr[5]~q ),
	.m_addr_6(\sdram|m_addr[6]~q ),
	.m_addr_7(\sdram|m_addr[7]~q ),
	.m_addr_8(\sdram|m_addr[8]~q ),
	.m_addr_9(\sdram|m_addr[9]~q ),
	.oe1(\sdram|oe~q ),
	.m_addr_10(\sdram|m_addr[10]~q ),
	.m_addr_11(\sdram|m_addr[11]~q ),
	.m_addr_12(\sdram|m_addr[12]~q ),
	.m_bank_0(\sdram|m_bank[0]~q ),
	.m_bank_1(\sdram|m_bank[1]~q ),
	.m_cmd_1(\sdram|m_cmd[1]~q ),
	.m_cmd_3(\sdram|m_cmd[3]~q ),
	.m_dqm_0(\sdram|m_dqm[0]~q ),
	.m_dqm_1(\sdram|m_dqm[1]~q ),
	.m_dqm_2(\sdram|m_dqm[2]~q ),
	.m_dqm_3(\sdram|m_dqm[3]~q ),
	.m_cmd_2(\sdram|m_cmd[2]~q ),
	.m_cmd_0(\sdram|m_cmd[0]~q ),
	.entries_1(\sdram|the_final_project_soc_sdram_input_efifo_module|entries[1]~q ),
	.entries_0(\sdram|the_final_project_soc_sdram_input_efifo_module|entries[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.last_cycle(\mm_interconnect_0|cmd_mux_006|last_cycle~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_006|saved_grant[1]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_006|WideOr1~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_006|src_payload~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux_006|src_data[68]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_006|src_data[48]~combout ),
	.src_data_62(\mm_interconnect_0|cmd_mux_006|src_data[62]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_006|src_data[49]~combout ),
	.src_data_51(\mm_interconnect_0|cmd_mux_006|src_data[51]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_006|src_data[50]~combout ),
	.src_data_53(\mm_interconnect_0|cmd_mux_006|src_data[53]~combout ),
	.src_data_52(\mm_interconnect_0|cmd_mux_006|src_data[52]~combout ),
	.src_data_55(\mm_interconnect_0|cmd_mux_006|src_data[55]~combout ),
	.src_data_54(\mm_interconnect_0|cmd_mux_006|src_data[54]~combout ),
	.src_data_57(\mm_interconnect_0|cmd_mux_006|src_data[57]~combout ),
	.src_data_56(\mm_interconnect_0|cmd_mux_006|src_data[56]~combout ),
	.src_data_59(\mm_interconnect_0|cmd_mux_006|src_data[59]~combout ),
	.src_data_58(\mm_interconnect_0|cmd_mux_006|src_data[58]~combout ),
	.src_data_61(\mm_interconnect_0|cmd_mux_006|src_data[61]~combout ),
	.src_data_60(\mm_interconnect_0|cmd_mux_006|src_data[60]~combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_006|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_006|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_006|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_006|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_006|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_006|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_006|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_006|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_006|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_006|src_data[47]~combout ),
	.out_data_buffer_32(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_321(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[32]~q ),
	.out_data_buffer_33(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_331(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[33]~q ),
	.out_data_buffer_34(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_341(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[34]~q ),
	.out_data_buffer_35(\mm_interconnect_0|crosser_001|clock_xer|out_data_buffer[35]~q ),
	.out_data_buffer_351(\mm_interconnect_0|crosser_003|clock_xer|out_data_buffer[35]~q ),
	.m_data_0(\sdram|m_data[0]~q ),
	.m_data_1(\sdram|m_data[1]~q ),
	.m_data_2(\sdram|m_data[2]~q ),
	.m_data_3(\sdram|m_data[3]~q ),
	.m_data_4(\sdram|m_data[4]~q ),
	.m_data_5(\sdram|m_data[5]~q ),
	.m_data_6(\sdram|m_data[6]~q ),
	.m_data_7(\sdram|m_data[7]~q ),
	.m_data_8(\sdram|m_data[8]~q ),
	.m_data_9(\sdram|m_data[9]~q ),
	.m_data_10(\sdram|m_data[10]~q ),
	.m_data_11(\sdram|m_data[11]~q ),
	.m_data_12(\sdram|m_data[12]~q ),
	.m_data_13(\sdram|m_data[13]~q ),
	.m_data_14(\sdram|m_data[14]~q ),
	.m_data_15(\sdram|m_data[15]~q ),
	.m_data_16(\sdram|m_data[16]~q ),
	.m_data_17(\sdram|m_data[17]~q ),
	.m_data_18(\sdram|m_data[18]~q ),
	.m_data_19(\sdram|m_data[19]~q ),
	.m_data_20(\sdram|m_data[20]~q ),
	.m_data_21(\sdram|m_data[21]~q ),
	.m_data_22(\sdram|m_data[22]~q ),
	.m_data_23(\sdram|m_data[23]~q ),
	.m_data_24(\sdram|m_data[24]~q ),
	.m_data_25(\sdram|m_data[25]~q ),
	.m_data_26(\sdram|m_data[26]~q ),
	.m_data_27(\sdram|m_data[27]~q ),
	.m_data_28(\sdram|m_data[28]~q ),
	.m_data_29(\sdram|m_data[29]~q ),
	.m_data_30(\sdram|m_data[30]~q ),
	.m_data_31(\sdram|m_data[31]~q ),
	.src_payload1(\mm_interconnect_0|cmd_mux_006|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_006|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_006|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_006|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_006|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_006|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_006|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_006|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_006|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_006|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_006|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_006|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_006|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_006|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_006|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_006|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_006|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_006|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_006|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_006|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_006|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_006|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_006|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_006|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_006|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_006|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_006|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_006|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_006|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_006|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_006|src_payload~31_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_006|src_payload~32_combout ),
	.za_valid1(\sdram|za_valid~q ),
	.za_data_0(\sdram|za_data[0]~q ),
	.za_data_1(\sdram|za_data[1]~q ),
	.za_data_2(\sdram|za_data[2]~q ),
	.za_data_3(\sdram|za_data[3]~q ),
	.za_data_4(\sdram|za_data[4]~q ),
	.za_data_11(\sdram|za_data[11]~q ),
	.za_data_13(\sdram|za_data[13]~q ),
	.za_data_16(\sdram|za_data[16]~q ),
	.za_data_12(\sdram|za_data[12]~q ),
	.za_data_5(\sdram|za_data[5]~q ),
	.za_data_14(\sdram|za_data[14]~q ),
	.za_data_15(\sdram|za_data[15]~q ),
	.za_data_21(\sdram|za_data[21]~q ),
	.za_data_18(\sdram|za_data[18]~q ),
	.za_data_17(\sdram|za_data[17]~q ),
	.za_data_31(\sdram|za_data[31]~q ),
	.za_data_30(\sdram|za_data[30]~q ),
	.za_data_29(\sdram|za_data[29]~q ),
	.za_data_28(\sdram|za_data[28]~q ),
	.za_data_27(\sdram|za_data[27]~q ),
	.za_data_26(\sdram|za_data[26]~q ),
	.za_data_25(\sdram|za_data[25]~q ),
	.za_data_10(\sdram|za_data[10]~q ),
	.za_data_24(\sdram|za_data[24]~q ),
	.za_data_9(\sdram|za_data[9]~q ),
	.za_data_23(\sdram|za_data[23]~q ),
	.za_data_8(\sdram|za_data[8]~q ),
	.za_data_22(\sdram|za_data[22]~q ),
	.za_data_7(\sdram|za_data[7]~q ),
	.za_data_6(\sdram|za_data[6]~q ),
	.za_data_20(\sdram|za_data[20]~q ),
	.za_data_19(\sdram|za_data[19]~q ),
	.m0_write(\mm_interconnect_0|sdram_s1_agent|m0_write~2_combout ),
	.sdram_wire_dq_0(\sdram_wire_dq[0]~input_o ),
	.sdram_wire_dq_1(\sdram_wire_dq[1]~input_o ),
	.sdram_wire_dq_2(\sdram_wire_dq[2]~input_o ),
	.sdram_wire_dq_3(\sdram_wire_dq[3]~input_o ),
	.sdram_wire_dq_4(\sdram_wire_dq[4]~input_o ),
	.sdram_wire_dq_5(\sdram_wire_dq[5]~input_o ),
	.sdram_wire_dq_6(\sdram_wire_dq[6]~input_o ),
	.sdram_wire_dq_7(\sdram_wire_dq[7]~input_o ),
	.sdram_wire_dq_8(\sdram_wire_dq[8]~input_o ),
	.sdram_wire_dq_9(\sdram_wire_dq[9]~input_o ),
	.sdram_wire_dq_10(\sdram_wire_dq[10]~input_o ),
	.sdram_wire_dq_11(\sdram_wire_dq[11]~input_o ),
	.sdram_wire_dq_12(\sdram_wire_dq[12]~input_o ),
	.sdram_wire_dq_13(\sdram_wire_dq[13]~input_o ),
	.sdram_wire_dq_14(\sdram_wire_dq[14]~input_o ),
	.sdram_wire_dq_15(\sdram_wire_dq[15]~input_o ),
	.sdram_wire_dq_16(\sdram_wire_dq[16]~input_o ),
	.sdram_wire_dq_17(\sdram_wire_dq[17]~input_o ),
	.sdram_wire_dq_18(\sdram_wire_dq[18]~input_o ),
	.sdram_wire_dq_19(\sdram_wire_dq[19]~input_o ),
	.sdram_wire_dq_20(\sdram_wire_dq[20]~input_o ),
	.sdram_wire_dq_21(\sdram_wire_dq[21]~input_o ),
	.sdram_wire_dq_22(\sdram_wire_dq[22]~input_o ),
	.sdram_wire_dq_23(\sdram_wire_dq[23]~input_o ),
	.sdram_wire_dq_24(\sdram_wire_dq[24]~input_o ),
	.sdram_wire_dq_25(\sdram_wire_dq[25]~input_o ),
	.sdram_wire_dq_26(\sdram_wire_dq[26]~input_o ),
	.sdram_wire_dq_27(\sdram_wire_dq[27]~input_o ),
	.sdram_wire_dq_28(\sdram_wire_dq[28]~input_o ),
	.sdram_wire_dq_29(\sdram_wire_dq[29]~input_o ),
	.sdram_wire_dq_30(\sdram_wire_dq[30]~input_o ),
	.sdram_wire_dq_31(\sdram_wire_dq[31]~input_o ));

final_project_soc_final_project_soc_onchip_memory2_0 onchip_memory2_0(
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.uav_write(\mm_interconnect_0|nios2_qsys_0_data_master_translator|uav_write~0_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_009|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr1(\mm_interconnect_0|cmd_mux_009|WideOr1~combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_009|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_009|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_009|src_data[39]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_009|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_009|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_009|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_009|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_009|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_009|src_payload~5_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_009|src_data[33]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_009|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_009|src_payload~7_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_009|src_data[34]~combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_009|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_009|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_009|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_009|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_009|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_009|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_009|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_009|src_payload~15_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_009|src_data[35]~combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_009|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_009|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_009|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_009|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_009|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_009|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_009|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_009|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_009|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_009|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_009|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_009|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_009|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_009|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_009|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_009|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

final_project_soc_final_project_soc_audio audio(
	.clk_0(\audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|clk[0] ),
	.readdata_0(\audio|readdata[0]~q ),
	.readdata_1(\audio|readdata[1]~q ),
	.readdata_2(\audio|readdata[2]~q ),
	.readdata_3(\audio|readdata[3]~q ),
	.readdata_4(\audio|readdata[4]~q ),
	.readdata_11(\audio|readdata[11]~q ),
	.readdata_13(\audio|readdata[13]~q ),
	.readdata_16(\audio|readdata[16]~q ),
	.readdata_12(\audio|readdata[12]~q ),
	.readdata_5(\audio|readdata[5]~q ),
	.readdata_14(\audio|readdata[14]~q ),
	.readdata_15(\audio|readdata[15]~q ),
	.readdata_21(\audio|readdata[21]~q ),
	.readdata_18(\audio|readdata[18]~q ),
	.readdata_17(\audio|readdata[17]~q ),
	.readdata_31(\audio|readdata[31]~q ),
	.readdata_30(\audio|readdata[30]~q ),
	.readdata_29(\audio|readdata[29]~q ),
	.readdata_28(\audio|readdata[28]~q ),
	.readdata_27(\audio|readdata[27]~q ),
	.readdata_26(\audio|readdata[26]~q ),
	.readdata_25(\audio|readdata[25]~q ),
	.readdata_10(\audio|readdata[10]~q ),
	.readdata_24(\audio|readdata[24]~q ),
	.readdata_9(\audio|readdata[9]~q ),
	.readdata_23(\audio|readdata[23]~q ),
	.readdata_8(\audio|readdata[8]~q ),
	.readdata_22(\audio|readdata[22]~q ),
	.readdata_7(\audio|readdata[7]~q ),
	.readdata_6(\audio|readdata[6]~q ),
	.readdata_20(\audio|readdata[20]~q ),
	.readdata_19(\audio|readdata[19]~q ),
	.irq1(\audio|irq~q ),
	.serial_audio_out_data(\audio|Audio_Out_Serializer|serial_audio_out_data~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux|saved_grant[0]~q ),
	.out_data_buffer_3(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[3]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux|src_data[39]~combout ),
	.WideOr1(\mm_interconnect_0|cmd_mux|WideOr1~combout ),
	.mem_used_1(\mm_interconnect_0|audio_avalon_audio_slave_agent_rsp_fifo|mem_used[1]~q ),
	.last_cycle(\mm_interconnect_0|cmd_mux|last_cycle~0_combout ),
	.nonposted_write_endofpacket(\mm_interconnect_0|audio_avalon_audio_slave_agent|nonposted_write_endofpacket~0_combout ),
	.src_payload(\mm_interconnect_0|cmd_mux|src_payload~0_combout ),
	.src_data_68(\mm_interconnect_0|cmd_mux|src_data[68]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux|src_payload~3_combout ),
	.out_data_buffer_0(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\mm_interconnect_0|crosser|clock_xer|out_data_buffer[2]~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux|src_payload~31_combout ),
	.GND_port(\~GND~combout ),
	.audio_wire_DACLRCK(\audio_wire_DACLRCK~input_o ),
	.audio_wire_BCLK(\audio_wire_BCLK~input_o ),
	.audio_wire_ADCLRCK(\audio_wire_ADCLRCK~input_o ),
	.audio_wire_ADCDAT(\audio_wire_ADCDAT~input_o ));

final_project_soc_altera_reset_controller_2 rst_controller_002(
	.wire_pll7_clk_0(\sdram_pll|sd1|wire_pll7_clk[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.reset_reset_n(\reset_reset_n~input_o ));

final_project_soc_altera_reset_controller_1 rst_controller_001(
	.locked(\audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|locked ),
	.clk_0(\audio_pll_0|audio_pll|PLL_for_DE_Series_Boards|auto_generated|clk[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

final_project_soc_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

final_project_soc_altera_irq_clock_crosser irq_synchronizer(
	.irq(\audio|irq~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.dreg_1(\irq_synchronizer|sync|sync[0].u|dreg[1]~q ),
	.clk_clk(\clk_clk~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~4_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .lut_mask = 16'h8BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .sum_lutc_input = "datac";

assign \audio_config_wire_SDAT~input_o  = audio_config_wire_SDAT;

assign \sdram_wire_dq[0]~input_o  = sdram_wire_dq[0];

assign \sdram_wire_dq[1]~input_o  = sdram_wire_dq[1];

assign \sdram_wire_dq[2]~input_o  = sdram_wire_dq[2];

assign \sdram_wire_dq[3]~input_o  = sdram_wire_dq[3];

assign \sdram_wire_dq[4]~input_o  = sdram_wire_dq[4];

assign \sdram_wire_dq[5]~input_o  = sdram_wire_dq[5];

assign \sdram_wire_dq[6]~input_o  = sdram_wire_dq[6];

assign \sdram_wire_dq[7]~input_o  = sdram_wire_dq[7];

assign \sdram_wire_dq[8]~input_o  = sdram_wire_dq[8];

assign \sdram_wire_dq[9]~input_o  = sdram_wire_dq[9];

assign \sdram_wire_dq[10]~input_o  = sdram_wire_dq[10];

assign \sdram_wire_dq[11]~input_o  = sdram_wire_dq[11];

assign \sdram_wire_dq[12]~input_o  = sdram_wire_dq[12];

assign \sdram_wire_dq[13]~input_o  = sdram_wire_dq[13];

assign \sdram_wire_dq[14]~input_o  = sdram_wire_dq[14];

assign \sdram_wire_dq[15]~input_o  = sdram_wire_dq[15];

assign \sdram_wire_dq[16]~input_o  = sdram_wire_dq[16];

assign \sdram_wire_dq[17]~input_o  = sdram_wire_dq[17];

assign \sdram_wire_dq[18]~input_o  = sdram_wire_dq[18];

assign \sdram_wire_dq[19]~input_o  = sdram_wire_dq[19];

assign \sdram_wire_dq[20]~input_o  = sdram_wire_dq[20];

assign \sdram_wire_dq[21]~input_o  = sdram_wire_dq[21];

assign \sdram_wire_dq[22]~input_o  = sdram_wire_dq[22];

assign \sdram_wire_dq[23]~input_o  = sdram_wire_dq[23];

assign \sdram_wire_dq[24]~input_o  = sdram_wire_dq[24];

assign \sdram_wire_dq[25]~input_o  = sdram_wire_dq[25];

assign \sdram_wire_dq[26]~input_o  = sdram_wire_dq[26];

assign \sdram_wire_dq[27]~input_o  = sdram_wire_dq[27];

assign \sdram_wire_dq[28]~input_o  = sdram_wire_dq[28];

assign \sdram_wire_dq[29]~input_o  = sdram_wire_dq[29];

assign \sdram_wire_dq[30]~input_o  = sdram_wire_dq[30];

assign \sdram_wire_dq[31]~input_o  = sdram_wire_dq[31];

assign \clk_clk~input_o  = clk_clk;

assign \unused_sdram_areset_conduit_export~input_o  = unused_sdram_areset_conduit_export;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \audio_wire_DACLRCK~input_o  = audio_wire_DACLRCK;

assign \audio_wire_BCLK~input_o  = audio_wire_BCLK;

assign \audio_wire_ADCLRCK~input_o  = audio_wire_ADCLRCK;

assign \audio_wire_ADCDAT~input_o  = audio_wire_ADCDAT;

assign audio_config_wire_SCLK = \audio_config|Serial_Bus_Controller|serial_clk~0_combout ;

assign audio_wire_DACDAT = \audio|Audio_Out_Serializer|serial_audio_out_data~q ;

assign ledg_wire_export[0] = \ledg|data_out[0]~q ;

assign ledg_wire_export[1] = \ledg|data_out[1]~q ;

assign ledg_wire_export[2] = \ledg|data_out[2]~q ;

assign ledg_wire_export[3] = \ledg|data_out[3]~q ;

assign ledg_wire_export[4] = \ledg|data_out[4]~q ;

assign ledg_wire_export[5] = \ledg|data_out[5]~q ;

assign ledg_wire_export[6] = \ledg|data_out[6]~q ;

assign ledg_wire_export[7] = \ledg|data_out[7]~q ;

assign ledr_wire_export[0] = \ledr|data_out[0]~q ;

assign ledr_wire_export[1] = \ledr|data_out[1]~q ;

assign ledr_wire_export[2] = \ledr|data_out[2]~q ;

assign ledr_wire_export[3] = \ledr|data_out[3]~q ;

assign ledr_wire_export[4] = \ledr|data_out[4]~q ;

assign ledr_wire_export[5] = \ledr|data_out[5]~q ;

assign ledr_wire_export[6] = \ledr|data_out[6]~q ;

assign ledr_wire_export[7] = \ledr|data_out[7]~q ;

assign ledr_wire_export[8] = \ledr|data_out[8]~q ;

assign ledr_wire_export[9] = \ledr|data_out[9]~q ;

assign ledr_wire_export[10] = \ledr|data_out[10]~q ;

assign ledr_wire_export[11] = \ledr|data_out[11]~q ;

assign ledr_wire_export[12] = \ledr|data_out[12]~q ;

assign ledr_wire_export[13] = \ledr|data_out[13]~q ;

assign ledr_wire_export[14] = \ledr|data_out[14]~q ;

assign ledr_wire_export[15] = \ledr|data_out[15]~q ;

assign ledr_wire_export[16] = \ledr|data_out[16]~q ;

assign ledr_wire_export[17] = \ledr|data_out[17]~q ;

assign sdram_clk_clk = \sdram_pll|sd1|wire_pll7_clk[1] ;

assign sdram_wire_addr[0] = \sdram|m_addr[0]~q ;

assign sdram_wire_addr[1] = \sdram|m_addr[1]~q ;

assign sdram_wire_addr[2] = \sdram|m_addr[2]~q ;

assign sdram_wire_addr[3] = \sdram|m_addr[3]~q ;

assign sdram_wire_addr[4] = \sdram|m_addr[4]~q ;

assign sdram_wire_addr[5] = \sdram|m_addr[5]~q ;

assign sdram_wire_addr[6] = \sdram|m_addr[6]~q ;

assign sdram_wire_addr[7] = \sdram|m_addr[7]~q ;

assign sdram_wire_addr[8] = \sdram|m_addr[8]~q ;

assign sdram_wire_addr[9] = \sdram|m_addr[9]~q ;

assign sdram_wire_addr[10] = \sdram|m_addr[10]~q ;

assign sdram_wire_addr[11] = \sdram|m_addr[11]~q ;

assign sdram_wire_addr[12] = \sdram|m_addr[12]~q ;

assign sdram_wire_ba[0] = \sdram|m_bank[0]~q ;

assign sdram_wire_ba[1] = \sdram|m_bank[1]~q ;

assign sdram_wire_cas_n = ~ \sdram|m_cmd[1]~q ;

assign sdram_wire_cke = vcc;

assign sdram_wire_cs_n = ~ \sdram|m_cmd[3]~q ;

assign sdram_wire_dqm[0] = \sdram|m_dqm[0]~q ;

assign sdram_wire_dqm[1] = \sdram|m_dqm[1]~q ;

assign sdram_wire_dqm[2] = \sdram|m_dqm[2]~q ;

assign sdram_wire_dqm[3] = \sdram|m_dqm[3]~q ;

assign sdram_wire_ras_n = ~ \sdram|m_cmd[2]~q ;

assign sdram_wire_we_n = ~ \sdram|m_cmd[0]~q ;

assign unused_sdram_locked_conduit_export = \sdram_pll|sd1|locked~combout ;

assign unused_sdram_phasedone_conduit_export = gnd;

cycloneive_io_obuf \audio_config_wire_SDAT~output (
	.i(\audio_config|Serial_Bus_Controller|serial_data~1_combout ),
	.oe(\audio_config|Serial_Bus_Controller|serial_data~2_combout ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(audio_config_wire_SDAT),
	.obar());
defparam \audio_config_wire_SDAT~output .bus_hold = "false";
defparam \audio_config_wire_SDAT~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[0]~output (
	.i(\sdram|m_data[0]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[0]),
	.obar());
defparam \sdram_wire_dq[0]~output .bus_hold = "false";
defparam \sdram_wire_dq[0]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[1]~output (
	.i(\sdram|m_data[1]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[1]),
	.obar());
defparam \sdram_wire_dq[1]~output .bus_hold = "false";
defparam \sdram_wire_dq[1]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[2]~output (
	.i(\sdram|m_data[2]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[2]),
	.obar());
defparam \sdram_wire_dq[2]~output .bus_hold = "false";
defparam \sdram_wire_dq[2]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[3]~output (
	.i(\sdram|m_data[3]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[3]),
	.obar());
defparam \sdram_wire_dq[3]~output .bus_hold = "false";
defparam \sdram_wire_dq[3]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[4]~output (
	.i(\sdram|m_data[4]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[4]),
	.obar());
defparam \sdram_wire_dq[4]~output .bus_hold = "false";
defparam \sdram_wire_dq[4]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[5]~output (
	.i(\sdram|m_data[5]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[5]),
	.obar());
defparam \sdram_wire_dq[5]~output .bus_hold = "false";
defparam \sdram_wire_dq[5]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[6]~output (
	.i(\sdram|m_data[6]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[6]),
	.obar());
defparam \sdram_wire_dq[6]~output .bus_hold = "false";
defparam \sdram_wire_dq[6]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[7]~output (
	.i(\sdram|m_data[7]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[7]),
	.obar());
defparam \sdram_wire_dq[7]~output .bus_hold = "false";
defparam \sdram_wire_dq[7]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[8]~output (
	.i(\sdram|m_data[8]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[8]),
	.obar());
defparam \sdram_wire_dq[8]~output .bus_hold = "false";
defparam \sdram_wire_dq[8]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[9]~output (
	.i(\sdram|m_data[9]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[9]),
	.obar());
defparam \sdram_wire_dq[9]~output .bus_hold = "false";
defparam \sdram_wire_dq[9]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[10]~output (
	.i(\sdram|m_data[10]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[10]),
	.obar());
defparam \sdram_wire_dq[10]~output .bus_hold = "false";
defparam \sdram_wire_dq[10]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[11]~output (
	.i(\sdram|m_data[11]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[11]),
	.obar());
defparam \sdram_wire_dq[11]~output .bus_hold = "false";
defparam \sdram_wire_dq[11]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[12]~output (
	.i(\sdram|m_data[12]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[12]),
	.obar());
defparam \sdram_wire_dq[12]~output .bus_hold = "false";
defparam \sdram_wire_dq[12]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[13]~output (
	.i(\sdram|m_data[13]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[13]),
	.obar());
defparam \sdram_wire_dq[13]~output .bus_hold = "false";
defparam \sdram_wire_dq[13]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[14]~output (
	.i(\sdram|m_data[14]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[14]),
	.obar());
defparam \sdram_wire_dq[14]~output .bus_hold = "false";
defparam \sdram_wire_dq[14]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[15]~output (
	.i(\sdram|m_data[15]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[15]),
	.obar());
defparam \sdram_wire_dq[15]~output .bus_hold = "false";
defparam \sdram_wire_dq[15]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[16]~output (
	.i(\sdram|m_data[16]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[16]),
	.obar());
defparam \sdram_wire_dq[16]~output .bus_hold = "false";
defparam \sdram_wire_dq[16]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[17]~output (
	.i(\sdram|m_data[17]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[17]),
	.obar());
defparam \sdram_wire_dq[17]~output .bus_hold = "false";
defparam \sdram_wire_dq[17]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[18]~output (
	.i(\sdram|m_data[18]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[18]),
	.obar());
defparam \sdram_wire_dq[18]~output .bus_hold = "false";
defparam \sdram_wire_dq[18]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[19]~output (
	.i(\sdram|m_data[19]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[19]),
	.obar());
defparam \sdram_wire_dq[19]~output .bus_hold = "false";
defparam \sdram_wire_dq[19]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[20]~output (
	.i(\sdram|m_data[20]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[20]),
	.obar());
defparam \sdram_wire_dq[20]~output .bus_hold = "false";
defparam \sdram_wire_dq[20]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[21]~output (
	.i(\sdram|m_data[21]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[21]),
	.obar());
defparam \sdram_wire_dq[21]~output .bus_hold = "false";
defparam \sdram_wire_dq[21]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[22]~output (
	.i(\sdram|m_data[22]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[22]),
	.obar());
defparam \sdram_wire_dq[22]~output .bus_hold = "false";
defparam \sdram_wire_dq[22]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[23]~output (
	.i(\sdram|m_data[23]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[23]),
	.obar());
defparam \sdram_wire_dq[23]~output .bus_hold = "false";
defparam \sdram_wire_dq[23]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[24]~output (
	.i(\sdram|m_data[24]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[24]),
	.obar());
defparam \sdram_wire_dq[24]~output .bus_hold = "false";
defparam \sdram_wire_dq[24]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[25]~output (
	.i(\sdram|m_data[25]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[25]),
	.obar());
defparam \sdram_wire_dq[25]~output .bus_hold = "false";
defparam \sdram_wire_dq[25]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[26]~output (
	.i(\sdram|m_data[26]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[26]),
	.obar());
defparam \sdram_wire_dq[26]~output .bus_hold = "false";
defparam \sdram_wire_dq[26]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[27]~output (
	.i(\sdram|m_data[27]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[27]),
	.obar());
defparam \sdram_wire_dq[27]~output .bus_hold = "false";
defparam \sdram_wire_dq[27]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[28]~output (
	.i(\sdram|m_data[28]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[28]),
	.obar());
defparam \sdram_wire_dq[28]~output .bus_hold = "false";
defparam \sdram_wire_dq[28]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[29]~output (
	.i(\sdram|m_data[29]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[29]),
	.obar());
defparam \sdram_wire_dq[29]~output .bus_hold = "false";
defparam \sdram_wire_dq[29]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[30]~output (
	.i(\sdram|m_data[30]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[30]),
	.obar());
defparam \sdram_wire_dq[30]~output .bus_hold = "false";
defparam \sdram_wire_dq[30]~output .open_drain_output = "false";

cycloneive_io_obuf \sdram_wire_dq[31]~output (
	.i(\sdram|m_data[31]~q ),
	.oe(\sdram|oe~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(sdram_wire_dq[31]),
	.obar());
defparam \sdram_wire_dq[31]~output .bus_hold = "false";
defparam \sdram_wire_dq[31]~output .open_drain_output = "false";

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0 (
	.dataa(\~GND~combout ),
	.datab(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 16'hBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .lut_mask = 16'h9696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~2_combout ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .lut_mask = 16'hBEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14 .lut_mask = 16'hDDF5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|ir_out[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal6~0_combout ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~11_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8 .lut_mask = 16'hFFDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|ir_out[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~9_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 .lut_mask = 16'hFFFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'h9696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 16'hFDFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'hFFBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'hFF7D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .lut_mask = 16'hBFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric_ident_writedata[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~15_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .lut_mask = 16'hFF6F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .lut_mask = 16'hFFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~19_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~20_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 (
	.dataa(\nios2_qsys_0|cpu|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\jtag_uart_0|final_project_soc_jtag_uart_0_alt_jtag_atlantic|tdo~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_irq_clock_crosser (
	irq,
	r_sync_rst,
	dreg_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	irq;
input 	r_sync_rst;
output 	dreg_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_std_synchronizer_bundle sync(
	.irq(irq),
	.r_sync_rst(r_sync_rst),
	.dreg_1(dreg_1),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_std_synchronizer_bundle (
	irq,
	r_sync_rst,
	dreg_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	irq;
input 	r_sync_rst;
output 	dreg_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_std_synchronizer \sync[0].u (
	.din(irq),
	.reset_n(r_sync_rst),
	.dreg_1(dreg_1),
	.clk(clk_clk));

endmodule

module final_project_soc_altera_std_synchronizer (
	din,
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module final_project_soc_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


final_project_soc_altera_reset_synchronizer_4 alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

final_project_soc_altera_reset_synchronizer_5 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 16'h5555;
defparam \altera_reset_synchronizer_int_chain[4]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.cout());
defparam \r_sync_rst_chain~1 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~1 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\altera_reset_synchronizer_int_chain[4]~q ),
	.datab(r_sync_rst1),
	.datac(gnd),
	.datad(\r_sync_rst_chain[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_reset_controller_1 (
	locked,
	clk_0,
	altera_reset_synchronizer_int_chain_out)/* synthesis synthesis_greybox=1 */;
input 	locked;
input 	clk_0;
output 	altera_reset_synchronizer_int_chain_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.locked(locked),
	.clk(clk_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out));

endmodule

module final_project_soc_altera_reset_synchronizer_1 (
	locked,
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=1 */;
input 	locked;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(locked),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(locked),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(locked),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module final_project_soc_altera_reset_controller_2 (
	wire_pll7_clk_0,
	altera_reset_synchronizer_int_chain_out,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.clk(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.reset_reset_n(reset_reset_n));

endmodule

module final_project_soc_altera_reset_synchronizer_3 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module final_project_soc_altera_reset_synchronizer_4 (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module final_project_soc_altera_reset_synchronizer_5 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_audio (
	clk_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_21,
	readdata_18,
	readdata_17,
	readdata_31,
	readdata_30,
	readdata_29,
	readdata_28,
	readdata_27,
	readdata_26,
	readdata_25,
	readdata_10,
	readdata_24,
	readdata_9,
	readdata_23,
	readdata_8,
	readdata_22,
	readdata_7,
	readdata_6,
	readdata_20,
	readdata_19,
	irq1,
	serial_audio_out_data,
	altera_reset_synchronizer_int_chain_out,
	saved_grant_0,
	out_data_buffer_3,
	src_data_38,
	src_data_39,
	WideOr1,
	mem_used_1,
	last_cycle,
	nonposted_write_endofpacket,
	src_payload,
	src_data_68,
	src_payload1,
	src_payload2,
	src_payload3,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	GND_port,
	audio_wire_DACLRCK,
	audio_wire_BCLK,
	audio_wire_ADCLRCK,
	audio_wire_ADCDAT)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_21;
output 	readdata_18;
output 	readdata_17;
output 	readdata_31;
output 	readdata_30;
output 	readdata_29;
output 	readdata_28;
output 	readdata_27;
output 	readdata_26;
output 	readdata_25;
output 	readdata_10;
output 	readdata_24;
output 	readdata_9;
output 	readdata_23;
output 	readdata_8;
output 	readdata_22;
output 	readdata_7;
output 	readdata_6;
output 	readdata_20;
output 	readdata_19;
output 	irq1;
output 	serial_audio_out_data;
input 	altera_reset_synchronizer_int_chain_out;
input 	saved_grant_0;
input 	out_data_buffer_3;
input 	src_data_38;
input 	src_data_39;
input 	WideOr1;
input 	mem_used_1;
input 	last_cycle;
input 	nonposted_write_endofpacket;
input 	src_payload;
input 	src_data_68;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	out_data_buffer_0;
input 	out_data_buffer_1;
input 	out_data_buffer_2;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	GND_port;
input 	audio_wire_DACLRCK;
input 	audio_wire_BCLK;
input 	audio_wire_ADCLRCK;
input 	audio_wire_ADCDAT;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \done_dac_channel_sync~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[0]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[5]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[2]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[1]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[7]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[6]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[5]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[4]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[3]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[2]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[1]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \Audio_Out_Serializer|left_channel_fifo_write_space[0]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[7]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[6]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[4]~q ;
wire \Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \Audio_Out_Serializer|right_channel_fifo_write_space[3]~q ;
wire \done_adc_channel_sync~q ;
wire \DAC_Left_Right_Clock_Edges|last_test_clk~q ;
wire \DAC_Left_Right_Clock_Edges|cur_test_clk~q ;
wire \comb~0_combout ;
wire \Bit_Clock_Edges|cur_test_clk~q ;
wire \Bit_Clock_Edges|last_test_clk~q ;
wire \Bit_Clock_Edges|falling_edge~combout ;
wire \done_dac_channel_sync~0_combout ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[0]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[1]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[2]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[3]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[4]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[3]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[5]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[4]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[5]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[6]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[7]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[2]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[1]~q ;
wire \Audio_In_Deserializer|left_audio_fifo_read_space[0]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[7]~q ;
wire \Audio_In_Deserializer|right_audio_fifo_read_space[6]~q ;
wire \ADC_Left_Right_Clock_Edges|last_test_clk~q ;
wire \ADC_Left_Right_Clock_Edges|cur_test_clk~q ;
wire \done_adc_channel_sync~0_combout ;
wire \comb~1_combout ;
wire \ADC_Left_Right_Clock_Edges|found_edge~combout ;
wire \read_interrupt_en~0_combout ;
wire \readdata[31]~26_combout ;
wire \clear_write_fifos~1_combout ;
wire \read_interrupt_en~q ;
wire \readdata~27_combout ;
wire \readdata~28_combout ;
wire \readdata[3]~29_combout ;
wire \write_interrupt_en~0_combout ;
wire \write_interrupt_en~q ;
wire \readdata~30_combout ;
wire \readdata~31_combout ;
wire \clear_read_fifos~0_combout ;
wire \clear_read_fifos~q ;
wire \readdata~32_combout ;
wire \readdata~33_combout ;
wire \clear_write_fifos~0_combout ;
wire \clear_write_fifos~q ;
wire \readdata~34_combout ;
wire \readdata~35_combout ;
wire \readdata[4]~0_combout ;
wire \readdata[31]~36_combout ;
wire \readdata[11]~9_combout ;
wire \readdata[13]~10_combout ;
wire \readdata[16]~11_combout ;
wire \readdata[12]~12_combout ;
wire \readdata[5]~6_combout ;
wire \readdata[14]~8_combout ;
wire \readdata[15]~7_combout ;
wire \readdata[21]~14_combout ;
wire \readdata[18]~13_combout ;
wire \readdata[17]~16_combout ;
wire \readdata[31]~15_combout ;
wire \readdata[30]~17_combout ;
wire \readdata[29]~18_combout ;
wire \readdata[28]~19_combout ;
wire \readdata[27]~20_combout ;
wire \readdata[26]~5_combout ;
wire \readdata[25]~4_combout ;
wire \readdata[10]~21_combout ;
wire \readdata[24]~3_combout ;
wire \write_interrupt~0_combout ;
wire \write_interrupt~1_combout ;
wire \write_interrupt~q ;
wire \readdata~37_combout ;
wire \readdata~38_combout ;
wire \readdata[23]~2_combout ;
wire \read_interrupt~0_combout ;
wire \read_interrupt~1_combout ;
wire \read_interrupt~q ;
wire \readdata~39_combout ;
wire \readdata~40_combout ;
wire \readdata[22]~1_combout ;
wire \readdata[7]~22_combout ;
wire \readdata[6]~24_combout ;
wire \readdata[20]~23_combout ;
wire \readdata[19]~25_combout ;
wire \irq~0_combout ;


final_project_soc_altera_up_audio_out_serializer Audio_Out_Serializer(
	.clk_0(clk_0),
	.done_dac_channel_sync(\done_dac_channel_sync~q ),
	.right_channel_fifo_write_space_0(\Audio_Out_Serializer|right_channel_fifo_write_space[0]~q ),
	.right_channel_fifo_write_space_5(\Audio_Out_Serializer|right_channel_fifo_write_space[5]~q ),
	.right_channel_fifo_write_space_2(\Audio_Out_Serializer|right_channel_fifo_write_space[2]~q ),
	.right_channel_fifo_write_space_1(\Audio_Out_Serializer|right_channel_fifo_write_space[1]~q ),
	.left_channel_fifo_write_space_7(\Audio_Out_Serializer|left_channel_fifo_write_space[7]~q ),
	.left_channel_fifo_write_space_6(\Audio_Out_Serializer|left_channel_fifo_write_space[6]~q ),
	.left_channel_fifo_write_space_5(\Audio_Out_Serializer|left_channel_fifo_write_space[5]~q ),
	.left_channel_fifo_write_space_4(\Audio_Out_Serializer|left_channel_fifo_write_space[4]~q ),
	.left_channel_fifo_write_space_3(\Audio_Out_Serializer|left_channel_fifo_write_space[3]~q ),
	.left_channel_fifo_write_space_2(\Audio_Out_Serializer|left_channel_fifo_write_space[2]~q ),
	.left_channel_fifo_write_space_1(\Audio_Out_Serializer|left_channel_fifo_write_space[1]~q ),
	.left_channel_fifo_write_space_0(\Audio_Out_Serializer|left_channel_fifo_write_space[0]~q ),
	.right_channel_fifo_write_space_7(\Audio_Out_Serializer|right_channel_fifo_write_space[7]~q ),
	.right_channel_fifo_write_space_6(\Audio_Out_Serializer|right_channel_fifo_write_space[6]~q ),
	.right_channel_fifo_write_space_4(\Audio_Out_Serializer|right_channel_fifo_write_space[4]~q ),
	.right_channel_fifo_write_space_3(\Audio_Out_Serializer|right_channel_fifo_write_space[3]~q ),
	.serial_audio_out_data1(serial_audio_out_data),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(\clear_write_fifos~q ),
	.last_test_clk(\DAC_Left_Right_Clock_Edges|last_test_clk~q ),
	.cur_test_clk(\DAC_Left_Right_Clock_Edges|cur_test_clk~q ),
	.comb(\comb~0_combout ),
	.falling_edge(\Bit_Clock_Edges|falling_edge~combout ),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.WideOr1(WideOr1),
	.mem_used_1(mem_used_1),
	.nonposted_write_endofpacket(nonposted_write_endofpacket),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.GND_port(GND_port));

final_project_soc_altera_up_audio_in_deserializer Audio_In_Deserializer(
	.clk_0(clk_0),
	.q_b_0(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_01(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_11(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_21(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_31(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_41(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_111(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_112(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_13(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_131(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_16(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_161(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_12(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_121(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_5(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_51(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_14(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_141(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_15(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_151(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_211(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_212(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_18(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_181(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_17(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_171(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_311(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_312(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_30(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_301(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_29(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_291(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_28(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_281(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_27(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_271(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_26(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_261(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_25(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_251(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_10(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_101(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_24(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_241(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_9(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_91(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_23(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_231(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_8(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_81(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_22(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_221(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_7(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_71(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_61(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_20(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_201(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_19(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_191(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.done_adc_channel_sync(\done_adc_channel_sync~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.cur_test_clk(\Bit_Clock_Edges|cur_test_clk~q ),
	.last_test_clk(\Bit_Clock_Edges|last_test_clk~q ),
	.falling_edge(\Bit_Clock_Edges|falling_edge~combout ),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.WideOr1(WideOr1),
	.mem_used_1(mem_used_1),
	.src_data_68(src_data_68),
	.right_audio_fifo_read_space_0(\Audio_In_Deserializer|right_audio_fifo_read_space[0]~q ),
	.right_audio_fifo_read_space_1(\Audio_In_Deserializer|right_audio_fifo_read_space[1]~q ),
	.right_audio_fifo_read_space_2(\Audio_In_Deserializer|right_audio_fifo_read_space[2]~q ),
	.clear_read_fifos(\clear_read_fifos~q ),
	.right_audio_fifo_read_space_3(\Audio_In_Deserializer|right_audio_fifo_read_space[3]~q ),
	.right_audio_fifo_read_space_4(\Audio_In_Deserializer|right_audio_fifo_read_space[4]~q ),
	.left_audio_fifo_read_space_3(\Audio_In_Deserializer|left_audio_fifo_read_space[3]~q ),
	.left_audio_fifo_read_space_5(\Audio_In_Deserializer|left_audio_fifo_read_space[5]~q ),
	.left_audio_fifo_read_space_4(\Audio_In_Deserializer|left_audio_fifo_read_space[4]~q ),
	.right_audio_fifo_read_space_5(\Audio_In_Deserializer|right_audio_fifo_read_space[5]~q ),
	.left_audio_fifo_read_space_6(\Audio_In_Deserializer|left_audio_fifo_read_space[6]~q ),
	.left_audio_fifo_read_space_7(\Audio_In_Deserializer|left_audio_fifo_read_space[7]~q ),
	.left_audio_fifo_read_space_2(\Audio_In_Deserializer|left_audio_fifo_read_space[2]~q ),
	.left_audio_fifo_read_space_1(\Audio_In_Deserializer|left_audio_fifo_read_space[1]~q ),
	.left_audio_fifo_read_space_0(\Audio_In_Deserializer|left_audio_fifo_read_space[0]~q ),
	.right_audio_fifo_read_space_7(\Audio_In_Deserializer|right_audio_fifo_read_space[7]~q ),
	.right_audio_fifo_read_space_6(\Audio_In_Deserializer|right_audio_fifo_read_space[6]~q ),
	.last_test_clk1(\ADC_Left_Right_Clock_Edges|last_test_clk~q ),
	.cur_test_clk1(\ADC_Left_Right_Clock_Edges|cur_test_clk~q ),
	.comb(\comb~1_combout ),
	.found_edge(\ADC_Left_Right_Clock_Edges|found_edge~combout ),
	.GND_port(GND_port),
	.audio_wire_ADCDAT(audio_wire_ADCDAT));

final_project_soc_altera_up_clock_edge_2 DAC_Left_Right_Clock_Edges(
	.clk(clk_0),
	.last_test_clk1(\DAC_Left_Right_Clock_Edges|last_test_clk~q ),
	.cur_test_clk1(\DAC_Left_Right_Clock_Edges|cur_test_clk~q ),
	.test_clk(audio_wire_DACLRCK));

final_project_soc_altera_up_clock_edge ADC_Left_Right_Clock_Edges(
	.clk(clk_0),
	.last_test_clk1(\ADC_Left_Right_Clock_Edges|last_test_clk~q ),
	.cur_test_clk1(\ADC_Left_Right_Clock_Edges|cur_test_clk~q ),
	.found_edge1(\ADC_Left_Right_Clock_Edges|found_edge~combout ),
	.test_clk(audio_wire_ADCLRCK));

final_project_soc_altera_up_clock_edge_1 Bit_Clock_Edges(
	.clk(clk_0),
	.cur_test_clk1(\Bit_Clock_Edges|cur_test_clk~q ),
	.last_test_clk1(\Bit_Clock_Edges|last_test_clk~q ),
	.falling_edge1(\Bit_Clock_Edges|falling_edge~combout ),
	.test_clk(audio_wire_BCLK));

dffeas done_dac_channel_sync(
	.clk(clk_0),
	.d(\done_dac_channel_sync~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\done_dac_channel_sync~q ),
	.prn(vcc));
defparam done_dac_channel_sync.is_wysiwyg = "true";
defparam done_dac_channel_sync.power_up = "low";

dffeas done_adc_channel_sync(
	.clk(clk_0),
	.d(\done_adc_channel_sync~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\done_adc_channel_sync~q ),
	.prn(vcc));
defparam done_adc_channel_sync.is_wysiwyg = "true";
defparam done_adc_channel_sync.power_up = "low";

cycloneive_lcell_comb \comb~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(gnd),
	.datad(\clear_write_fifos~q ),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hFF55;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \done_dac_channel_sync~0 (
	.dataa(\done_dac_channel_sync~q ),
	.datab(\DAC_Left_Right_Clock_Edges|last_test_clk~q ),
	.datac(gnd),
	.datad(\DAC_Left_Right_Clock_Edges|cur_test_clk~q ),
	.cin(gnd),
	.combout(\done_dac_channel_sync~0_combout ),
	.cout());
defparam \done_dac_channel_sync~0 .lut_mask = 16'hEEFF;
defparam \done_dac_channel_sync~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \done_adc_channel_sync~0 (
	.dataa(\done_adc_channel_sync~q ),
	.datab(\ADC_Left_Right_Clock_Edges|cur_test_clk~q ),
	.datac(gnd),
	.datad(\ADC_Left_Right_Clock_Edges|last_test_clk~q ),
	.cin(gnd),
	.combout(\done_adc_channel_sync~0_combout ),
	.cout());
defparam \done_adc_channel_sync~0 .lut_mask = 16'hEEFF;
defparam \done_adc_channel_sync~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(gnd),
	.datac(gnd),
	.datad(\clear_read_fifos~q ),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'hFF55;
defparam \comb~1 .sum_lutc_input = "datac";

dffeas \readdata[0] (
	.clk(clk_0),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_0),
	.d(\readdata~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_0),
	.d(\readdata~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_0),
	.d(\readdata~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_0),
	.d(\readdata[4]~0_combout ),
	.asdata(\Audio_In_Deserializer|right_audio_fifo_read_space[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_0),
	.d(\readdata[11]~9_combout ),
	.asdata(\Audio_In_Deserializer|left_audio_fifo_read_space[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_0),
	.d(\readdata[13]~10_combout ),
	.asdata(\Audio_In_Deserializer|left_audio_fifo_read_space[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_0),
	.d(\readdata[16]~11_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_0),
	.d(\readdata[12]~12_combout ),
	.asdata(\Audio_In_Deserializer|left_audio_fifo_read_space[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_0),
	.d(\readdata[5]~6_combout ),
	.asdata(\Audio_In_Deserializer|right_audio_fifo_read_space[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_0),
	.d(\readdata[14]~8_combout ),
	.asdata(\Audio_In_Deserializer|left_audio_fifo_read_space[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_0),
	.d(\readdata[15]~7_combout ),
	.asdata(\Audio_In_Deserializer|left_audio_fifo_read_space[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_0),
	.d(\readdata[21]~14_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_0),
	.d(\readdata[18]~13_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_0),
	.d(\readdata[17]~16_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_0),
	.d(\readdata[31]~15_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_0),
	.d(\readdata[30]~17_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_0),
	.d(\readdata[29]~18_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_0),
	.d(\readdata[28]~19_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_0),
	.d(\readdata[27]~20_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_0),
	.d(\readdata[26]~5_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_0),
	.d(\readdata[25]~4_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_0),
	.d(\readdata[10]~21_combout ),
	.asdata(\Audio_In_Deserializer|left_audio_fifo_read_space[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_0),
	.d(\readdata[24]~3_combout ),
	.asdata(\Audio_Out_Serializer|left_channel_fifo_write_space[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_0),
	.d(\readdata~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_0),
	.d(\readdata[23]~2_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_0),
	.d(\readdata~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_0),
	.d(\readdata[22]~1_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_0),
	.d(\readdata[7]~22_combout ),
	.asdata(\Audio_In_Deserializer|right_audio_fifo_read_space[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_0),
	.d(\readdata[6]~24_combout ),
	.asdata(\Audio_In_Deserializer|right_audio_fifo_read_space[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_0),
	.d(\readdata[20]~23_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_0),
	.d(\readdata[19]~25_combout ),
	.asdata(\Audio_Out_Serializer|right_channel_fifo_write_space[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\readdata[31]~36_combout ),
	.sload(src_data_39),
	.ena(\readdata[3]~29_combout ),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas irq(
	.clk(clk_0),
	.d(\irq~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(irq1),
	.prn(vcc));
defparam irq.is_wysiwyg = "true";
defparam irq.power_up = "low";

cycloneive_lcell_comb \read_interrupt_en~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(saved_grant_0),
	.datac(out_data_buffer_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_interrupt_en~0_combout ),
	.cout());
defparam \read_interrupt_en~0 .lut_mask = 16'hFEFE;
defparam \read_interrupt_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[31]~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\readdata[31]~26_combout ),
	.cout());
defparam \readdata[31]~26 .lut_mask = 16'hFF0F;
defparam \readdata[31]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \clear_write_fifos~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\readdata[31]~26_combout ),
	.datac(last_cycle),
	.datad(nonposted_write_endofpacket),
	.cin(gnd),
	.combout(\clear_write_fifos~1_combout ),
	.cout());
defparam \clear_write_fifos~1 .lut_mask = 16'hFFFD;
defparam \clear_write_fifos~1 .sum_lutc_input = "datac";

dffeas read_interrupt_en(
	.clk(clk_0),
	.d(\read_interrupt_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\clear_write_fifos~1_combout ),
	.q(\read_interrupt_en~q ),
	.prn(vcc));
defparam read_interrupt_en.is_wysiwyg = "true";
defparam read_interrupt_en.power_up = "low";

cycloneive_lcell_comb \readdata~27 (
	.dataa(src_data_39),
	.datab(\Audio_In_Deserializer|right_audio_fifo_read_space[0]~q ),
	.datac(src_data_38),
	.datad(\read_interrupt_en~q ),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hFFDE;
defparam \readdata~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~28 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(src_data_39),
	.datac(\readdata~27_combout ),
	.datad(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hFFBE;
defparam \readdata~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3]~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(nonposted_write_endofpacket),
	.datac(src_data_68),
	.datad(last_cycle),
	.cin(gnd),
	.combout(\readdata[3]~29_combout ),
	.cout());
defparam \readdata[3]~29 .lut_mask = 16'hFFFD;
defparam \readdata[3]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_interrupt_en~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(saved_grant_0),
	.datac(out_data_buffer_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_interrupt_en~0_combout ),
	.cout());
defparam \write_interrupt_en~0 .lut_mask = 16'hFEFE;
defparam \write_interrupt_en~0 .sum_lutc_input = "datac";

dffeas write_interrupt_en(
	.clk(clk_0),
	.d(\write_interrupt_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\clear_write_fifos~1_combout ),
	.q(\write_interrupt_en~q ),
	.prn(vcc));
defparam write_interrupt_en.is_wysiwyg = "true";
defparam write_interrupt_en.power_up = "low";

cycloneive_lcell_comb \readdata~30 (
	.dataa(src_data_38),
	.datab(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(src_data_39),
	.datad(\write_interrupt_en~q ),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hFFDE;
defparam \readdata~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~31 (
	.dataa(\Audio_In_Deserializer|right_audio_fifo_read_space[1]~q ),
	.datab(src_data_38),
	.datac(\readdata~30_combout ),
	.datad(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.cin(gnd),
	.combout(\readdata~31_combout ),
	.cout());
defparam \readdata~31 .lut_mask = 16'hFFBE;
defparam \readdata~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \clear_read_fifos~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(saved_grant_0),
	.datac(out_data_buffer_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\clear_read_fifos~0_combout ),
	.cout());
defparam \clear_read_fifos~0 .lut_mask = 16'hFEFE;
defparam \clear_read_fifos~0 .sum_lutc_input = "datac";

dffeas clear_read_fifos(
	.clk(clk_0),
	.d(\clear_read_fifos~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\clear_write_fifos~1_combout ),
	.q(\clear_read_fifos~q ),
	.prn(vcc));
defparam clear_read_fifos.is_wysiwyg = "true";
defparam clear_read_fifos.power_up = "low";

cycloneive_lcell_comb \readdata~32 (
	.dataa(src_data_39),
	.datab(\Audio_In_Deserializer|right_audio_fifo_read_space[2]~q ),
	.datac(src_data_38),
	.datad(\clear_read_fifos~q ),
	.cin(gnd),
	.combout(\readdata~32_combout ),
	.cout());
defparam \readdata~32 .lut_mask = 16'hFFDE;
defparam \readdata~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~33 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(src_data_39),
	.datac(\readdata~32_combout ),
	.datad(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.cin(gnd),
	.combout(\readdata~33_combout ),
	.cout());
defparam \readdata~33 .lut_mask = 16'hFFBE;
defparam \readdata~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \clear_write_fifos~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(saved_grant_0),
	.datac(out_data_buffer_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\clear_write_fifos~0_combout ),
	.cout());
defparam \clear_write_fifos~0 .lut_mask = 16'hFEFE;
defparam \clear_write_fifos~0 .sum_lutc_input = "datac";

dffeas clear_write_fifos(
	.clk(clk_0),
	.d(\clear_write_fifos~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\clear_write_fifos~1_combout ),
	.q(\clear_write_fifos~q ),
	.prn(vcc));
defparam clear_write_fifos.is_wysiwyg = "true";
defparam clear_write_fifos.power_up = "low";

cycloneive_lcell_comb \readdata~34 (
	.dataa(src_data_38),
	.datab(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(src_data_39),
	.datad(\clear_write_fifos~q ),
	.cin(gnd),
	.combout(\readdata~34_combout ),
	.cout());
defparam \readdata~34 .lut_mask = 16'hFFDE;
defparam \readdata~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~35 (
	.dataa(\Audio_In_Deserializer|right_audio_fifo_read_space[3]~q ),
	.datab(src_data_38),
	.datac(\readdata~34_combout ),
	.datad(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.cin(gnd),
	.combout(\readdata~35_combout ),
	.cout());
defparam \readdata~35 .lut_mask = 16'hFFBE;
defparam \readdata~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4]~0 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[4]~0_combout ),
	.cout());
defparam \readdata[4]~0 .lut_mask = 16'hAACC;
defparam \readdata[4]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[31]~36 (
	.dataa(gnd),
	.datab(src_data_38),
	.datac(src_data_39),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\readdata[31]~36_combout ),
	.cout());
defparam \readdata[31]~36 .lut_mask = 16'hF3FF;
defparam \readdata[31]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[11]~9 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[11]~9_combout ),
	.cout());
defparam \readdata[11]~9 .lut_mask = 16'hAACC;
defparam \readdata[11]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[13]~10 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[13]~10_combout ),
	.cout());
defparam \readdata[13]~10 .lut_mask = 16'hAACC;
defparam \readdata[13]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[16]~11 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[16]~11_combout ),
	.cout());
defparam \readdata[16]~11 .lut_mask = 16'hAACC;
defparam \readdata[16]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[12]~12 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[12]~12_combout ),
	.cout());
defparam \readdata[12]~12 .lut_mask = 16'hAACC;
defparam \readdata[12]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5]~6 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[5]~6_combout ),
	.cout());
defparam \readdata[5]~6 .lut_mask = 16'hAACC;
defparam \readdata[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[14]~8 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[14]~8_combout ),
	.cout());
defparam \readdata[14]~8 .lut_mask = 16'hAACC;
defparam \readdata[14]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[15]~7 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[15]~7_combout ),
	.cout());
defparam \readdata[15]~7 .lut_mask = 16'hAACC;
defparam \readdata[15]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[21]~14 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[21]~14_combout ),
	.cout());
defparam \readdata[21]~14 .lut_mask = 16'hAACC;
defparam \readdata[21]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[18]~13 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[18]~13_combout ),
	.cout());
defparam \readdata[18]~13 .lut_mask = 16'hAACC;
defparam \readdata[18]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[17]~16 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[17]~16_combout ),
	.cout());
defparam \readdata[17]~16 .lut_mask = 16'hAACC;
defparam \readdata[17]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[31]~15 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[31]~15_combout ),
	.cout());
defparam \readdata[31]~15 .lut_mask = 16'hAACC;
defparam \readdata[31]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[30]~17 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[30]~17_combout ),
	.cout());
defparam \readdata[30]~17 .lut_mask = 16'hAACC;
defparam \readdata[30]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[29]~18 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[29]~18_combout ),
	.cout());
defparam \readdata[29]~18 .lut_mask = 16'hAACC;
defparam \readdata[29]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[28]~19 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[28]~19_combout ),
	.cout());
defparam \readdata[28]~19 .lut_mask = 16'hAACC;
defparam \readdata[28]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[27]~20 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[27]~20_combout ),
	.cout());
defparam \readdata[27]~20 .lut_mask = 16'hAACC;
defparam \readdata[27]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[26]~5 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[26]~5_combout ),
	.cout());
defparam \readdata[26]~5 .lut_mask = 16'hAACC;
defparam \readdata[26]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[25]~4 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[25]~4_combout ),
	.cout());
defparam \readdata[25]~4 .lut_mask = 16'hAACC;
defparam \readdata[25]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[10]~21 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[10]~21_combout ),
	.cout());
defparam \readdata[10]~21 .lut_mask = 16'hAACC;
defparam \readdata[10]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[24]~3 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[24]~3_combout ),
	.cout());
defparam \readdata[24]~3 .lut_mask = 16'hAACC;
defparam \readdata[24]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_interrupt~0 (
	.dataa(\Audio_Out_Serializer|right_channel_fifo_write_space[5]~q ),
	.datab(\Audio_Out_Serializer|left_channel_fifo_write_space[6]~q ),
	.datac(\Audio_Out_Serializer|left_channel_fifo_write_space[5]~q ),
	.datad(\Audio_Out_Serializer|right_channel_fifo_write_space[6]~q ),
	.cin(gnd),
	.combout(\write_interrupt~0_combout ),
	.cout());
defparam \write_interrupt~0 .lut_mask = 16'hFFFE;
defparam \write_interrupt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_interrupt~1 (
	.dataa(\write_interrupt_en~q ),
	.datab(\Audio_Out_Serializer|left_channel_fifo_write_space[7]~q ),
	.datac(\Audio_Out_Serializer|right_channel_fifo_write_space[7]~q ),
	.datad(\write_interrupt~0_combout ),
	.cin(gnd),
	.combout(\write_interrupt~1_combout ),
	.cout());
defparam \write_interrupt~1 .lut_mask = 16'hFFFE;
defparam \write_interrupt~1 .sum_lutc_input = "datac";

dffeas write_interrupt(
	.clk(clk_0),
	.d(\write_interrupt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\write_interrupt~q ),
	.prn(vcc));
defparam write_interrupt.is_wysiwyg = "true";
defparam write_interrupt.power_up = "low";

cycloneive_lcell_comb \readdata~37 (
	.dataa(src_data_38),
	.datab(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(src_data_39),
	.datad(\write_interrupt~q ),
	.cin(gnd),
	.combout(\readdata~37_combout ),
	.cout());
defparam \readdata~37 .lut_mask = 16'hFFDE;
defparam \readdata~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~38 (
	.dataa(\Audio_In_Deserializer|left_audio_fifo_read_space[1]~q ),
	.datab(src_data_38),
	.datac(\readdata~37_combout ),
	.datad(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\readdata~38_combout ),
	.cout());
defparam \readdata~38 .lut_mask = 16'hFFBE;
defparam \readdata~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[23]~2 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[23]~2_combout ),
	.cout());
defparam \readdata[23]~2 .lut_mask = 16'hAACC;
defparam \readdata[23]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_interrupt~0 (
	.dataa(\Audio_In_Deserializer|right_audio_fifo_read_space[5]~q ),
	.datab(\Audio_In_Deserializer|left_audio_fifo_read_space[5]~q ),
	.datac(\Audio_In_Deserializer|left_audio_fifo_read_space[6]~q ),
	.datad(\Audio_In_Deserializer|right_audio_fifo_read_space[6]~q ),
	.cin(gnd),
	.combout(\read_interrupt~0_combout ),
	.cout());
defparam \read_interrupt~0 .lut_mask = 16'hFFFE;
defparam \read_interrupt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_interrupt~1 (
	.dataa(\read_interrupt_en~q ),
	.datab(\Audio_In_Deserializer|left_audio_fifo_read_space[7]~q ),
	.datac(\Audio_In_Deserializer|right_audio_fifo_read_space[7]~q ),
	.datad(\read_interrupt~0_combout ),
	.cin(gnd),
	.combout(\read_interrupt~1_combout ),
	.cout());
defparam \read_interrupt~1 .lut_mask = 16'hFFFE;
defparam \read_interrupt~1 .sum_lutc_input = "datac";

dffeas read_interrupt(
	.clk(clk_0),
	.d(\read_interrupt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!altera_reset_synchronizer_int_chain_out),
	.sload(gnd),
	.ena(vcc),
	.q(\read_interrupt~q ),
	.prn(vcc));
defparam read_interrupt.is_wysiwyg = "true";
defparam read_interrupt.power_up = "low";

cycloneive_lcell_comb \readdata~39 (
	.dataa(src_data_39),
	.datab(\Audio_In_Deserializer|left_audio_fifo_read_space[0]~q ),
	.datac(src_data_38),
	.datad(\read_interrupt~q ),
	.cin(gnd),
	.combout(\readdata~39_combout ),
	.cout());
defparam \readdata~39 .lut_mask = 16'hFFDE;
defparam \readdata~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~40 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(src_data_39),
	.datac(\readdata~39_combout ),
	.datad(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\readdata~40_combout ),
	.cout());
defparam \readdata~40 .lut_mask = 16'hFFBE;
defparam \readdata~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[22]~1 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[22]~1_combout ),
	.cout());
defparam \readdata[22]~1 .lut_mask = 16'hAACC;
defparam \readdata[22]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7]~22 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[7]~22_combout ),
	.cout());
defparam \readdata[7]~22 .lut_mask = 16'hAACC;
defparam \readdata[7]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6]~24 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[6]~24_combout ),
	.cout());
defparam \readdata[6]~24 .lut_mask = 16'hAACC;
defparam \readdata[6]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[20]~23 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[20]~23_combout ),
	.cout());
defparam \readdata[20]~23 .lut_mask = 16'hAACC;
defparam \readdata[20]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[19]~25 (
	.dataa(\Audio_In_Deserializer|Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datab(\Audio_In_Deserializer|Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata[19]~25_combout ),
	.cout());
defparam \readdata[19]~25 .lut_mask = 16'hAACC;
defparam \readdata[19]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \irq~0 (
	.dataa(\read_interrupt~q ),
	.datab(\write_interrupt~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\irq~0_combout ),
	.cout());
defparam \irq~0 .lut_mask = 16'hEEEE;
defparam \irq~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_audio_in_deserializer (
	clk_0,
	q_b_0,
	q_b_01,
	q_b_1,
	q_b_11,
	q_b_2,
	q_b_21,
	q_b_3,
	q_b_31,
	q_b_4,
	q_b_41,
	q_b_111,
	q_b_112,
	q_b_13,
	q_b_131,
	q_b_16,
	q_b_161,
	q_b_12,
	q_b_121,
	q_b_5,
	q_b_51,
	q_b_14,
	q_b_141,
	q_b_15,
	q_b_151,
	q_b_211,
	q_b_212,
	q_b_18,
	q_b_181,
	q_b_17,
	q_b_171,
	q_b_311,
	q_b_312,
	q_b_30,
	q_b_301,
	q_b_29,
	q_b_291,
	q_b_28,
	q_b_281,
	q_b_27,
	q_b_271,
	q_b_26,
	q_b_261,
	q_b_25,
	q_b_251,
	q_b_10,
	q_b_101,
	q_b_24,
	q_b_241,
	q_b_9,
	q_b_91,
	q_b_23,
	q_b_231,
	q_b_8,
	q_b_81,
	q_b_22,
	q_b_221,
	q_b_7,
	q_b_71,
	q_b_6,
	q_b_61,
	q_b_20,
	q_b_201,
	q_b_19,
	q_b_191,
	done_adc_channel_sync,
	altera_reset_synchronizer_int_chain_out,
	cur_test_clk,
	last_test_clk,
	falling_edge,
	src_data_38,
	src_data_39,
	WideOr1,
	mem_used_1,
	src_data_68,
	right_audio_fifo_read_space_0,
	right_audio_fifo_read_space_1,
	right_audio_fifo_read_space_2,
	clear_read_fifos,
	right_audio_fifo_read_space_3,
	right_audio_fifo_read_space_4,
	left_audio_fifo_read_space_3,
	left_audio_fifo_read_space_5,
	left_audio_fifo_read_space_4,
	right_audio_fifo_read_space_5,
	left_audio_fifo_read_space_6,
	left_audio_fifo_read_space_7,
	left_audio_fifo_read_space_2,
	left_audio_fifo_read_space_1,
	left_audio_fifo_read_space_0,
	right_audio_fifo_read_space_7,
	right_audio_fifo_read_space_6,
	last_test_clk1,
	cur_test_clk1,
	comb,
	found_edge,
	GND_port,
	audio_wire_ADCDAT)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
output 	q_b_0;
output 	q_b_01;
output 	q_b_1;
output 	q_b_11;
output 	q_b_2;
output 	q_b_21;
output 	q_b_3;
output 	q_b_31;
output 	q_b_4;
output 	q_b_41;
output 	q_b_111;
output 	q_b_112;
output 	q_b_13;
output 	q_b_131;
output 	q_b_16;
output 	q_b_161;
output 	q_b_12;
output 	q_b_121;
output 	q_b_5;
output 	q_b_51;
output 	q_b_14;
output 	q_b_141;
output 	q_b_15;
output 	q_b_151;
output 	q_b_211;
output 	q_b_212;
output 	q_b_18;
output 	q_b_181;
output 	q_b_17;
output 	q_b_171;
output 	q_b_311;
output 	q_b_312;
output 	q_b_30;
output 	q_b_301;
output 	q_b_29;
output 	q_b_291;
output 	q_b_28;
output 	q_b_281;
output 	q_b_27;
output 	q_b_271;
output 	q_b_26;
output 	q_b_261;
output 	q_b_25;
output 	q_b_251;
output 	q_b_10;
output 	q_b_101;
output 	q_b_24;
output 	q_b_241;
output 	q_b_9;
output 	q_b_91;
output 	q_b_23;
output 	q_b_231;
output 	q_b_8;
output 	q_b_81;
output 	q_b_22;
output 	q_b_221;
output 	q_b_7;
output 	q_b_71;
output 	q_b_6;
output 	q_b_61;
output 	q_b_20;
output 	q_b_201;
output 	q_b_19;
output 	q_b_191;
input 	done_adc_channel_sync;
input 	altera_reset_synchronizer_int_chain_out;
input 	cur_test_clk;
input 	last_test_clk;
input 	falling_edge;
input 	src_data_38;
input 	src_data_39;
input 	WideOr1;
input 	mem_used_1;
input 	src_data_68;
output 	right_audio_fifo_read_space_0;
output 	right_audio_fifo_read_space_1;
output 	right_audio_fifo_read_space_2;
input 	clear_read_fifos;
output 	right_audio_fifo_read_space_3;
output 	right_audio_fifo_read_space_4;
output 	left_audio_fifo_read_space_3;
output 	left_audio_fifo_read_space_5;
output 	left_audio_fifo_read_space_4;
output 	right_audio_fifo_read_space_5;
output 	left_audio_fifo_read_space_6;
output 	left_audio_fifo_read_space_7;
output 	left_audio_fifo_read_space_2;
output 	left_audio_fifo_read_space_1;
output 	left_audio_fifo_read_space_0;
output 	right_audio_fifo_read_space_7;
output 	right_audio_fifo_read_space_6;
input 	last_test_clk1;
input 	cur_test_clk1;
input 	comb;
input 	found_edge;
input 	GND_port;
input 	audio_wire_ADCDAT;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \Audio_Out_Bit_Counter|counting~q ;
wire \comb~0_combout ;
wire \data_in_shift_reg[0]~q ;
wire \comb~1_combout ;
wire \Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \comb~2_combout ;
wire \comb~3_combout ;
wire \Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \comb~4_combout ;
wire \data_in_shift_reg[1]~q ;
wire \data_in_shift_reg[2]~q ;
wire \data_in_shift_reg[3]~q ;
wire \data_in_shift_reg[4]~q ;
wire \data_in_shift_reg[11]~q ;
wire \data_in_shift_reg[13]~q ;
wire \data_in_shift_reg[16]~q ;
wire \data_in_shift_reg[12]~q ;
wire \data_in_shift_reg[5]~q ;
wire \data_in_shift_reg[14]~q ;
wire \data_in_shift_reg[15]~q ;
wire \data_in_shift_reg[21]~q ;
wire \data_in_shift_reg[18]~q ;
wire \data_in_shift_reg[17]~q ;
wire \data_in_shift_reg[31]~q ;
wire \data_in_shift_reg[30]~q ;
wire \data_in_shift_reg[29]~q ;
wire \data_in_shift_reg[28]~q ;
wire \data_in_shift_reg[27]~q ;
wire \data_in_shift_reg[26]~q ;
wire \data_in_shift_reg[25]~q ;
wire \data_in_shift_reg[10]~q ;
wire \data_in_shift_reg[24]~q ;
wire \data_in_shift_reg[9]~q ;
wire \data_in_shift_reg[23]~q ;
wire \data_in_shift_reg[8]~q ;
wire \data_in_shift_reg[22]~q ;
wire \data_in_shift_reg[7]~q ;
wire \data_in_shift_reg[6]~q ;
wire \data_in_shift_reg[20]~q ;
wire \data_in_shift_reg[19]~q ;
wire \data_in_shift_reg~0_combout ;
wire \data_in_shift_reg[9]~1_combout ;
wire \data_in_shift_reg~2_combout ;
wire \data_in_shift_reg~3_combout ;
wire \data_in_shift_reg~4_combout ;
wire \data_in_shift_reg~5_combout ;
wire \data_in_shift_reg~6_combout ;
wire \data_in_shift_reg~7_combout ;
wire \data_in_shift_reg~8_combout ;
wire \data_in_shift_reg~9_combout ;
wire \data_in_shift_reg~10_combout ;
wire \data_in_shift_reg~11_combout ;
wire \data_in_shift_reg~12_combout ;
wire \data_in_shift_reg~13_combout ;
wire \data_in_shift_reg~14_combout ;
wire \data_in_shift_reg~15_combout ;
wire \data_in_shift_reg~16_combout ;
wire \data_in_shift_reg~17_combout ;
wire \data_in_shift_reg~18_combout ;
wire \data_in_shift_reg~19_combout ;
wire \data_in_shift_reg~20_combout ;
wire \data_in_shift_reg~21_combout ;
wire \data_in_shift_reg~22_combout ;
wire \data_in_shift_reg~23_combout ;
wire \data_in_shift_reg~24_combout ;
wire \data_in_shift_reg~25_combout ;
wire \data_in_shift_reg~26_combout ;
wire \data_in_shift_reg~27_combout ;
wire \data_in_shift_reg~28_combout ;
wire \data_in_shift_reg~29_combout ;
wire \data_in_shift_reg~30_combout ;
wire \data_in_shift_reg~31_combout ;
wire \data_in_shift_reg~32_combout ;
wire \right_audio_fifo_read_space~0_combout ;
wire \right_audio_fifo_read_space~1_combout ;
wire \right_audio_fifo_read_space~2_combout ;
wire \right_audio_fifo_read_space~3_combout ;
wire \right_audio_fifo_read_space~4_combout ;
wire \left_audio_fifo_read_space~0_combout ;
wire \left_audio_fifo_read_space~1_combout ;
wire \left_audio_fifo_read_space~2_combout ;
wire \right_audio_fifo_read_space~5_combout ;
wire \left_audio_fifo_read_space~3_combout ;
wire \left_audio_fifo_read_space~4_combout ;
wire \left_audio_fifo_read_space~5_combout ;
wire \left_audio_fifo_read_space~6_combout ;
wire \left_audio_fifo_read_space~7_combout ;
wire \right_audio_fifo_read_space~6_combout ;
wire \right_audio_fifo_read_space~7_combout ;


final_project_soc_altera_up_sync_fifo_1 Audio_In_Right_Channel_FIFO(
	.clk_0(clk_0),
	.q_b_0(q_b_01),
	.q_b_1(q_b_11),
	.q_b_2(q_b_21),
	.q_b_3(q_b_31),
	.q_b_4(q_b_41),
	.q_b_11(q_b_112),
	.q_b_13(q_b_131),
	.q_b_16(q_b_161),
	.q_b_12(q_b_121),
	.q_b_5(q_b_51),
	.q_b_14(q_b_141),
	.q_b_15(q_b_151),
	.q_b_21(q_b_212),
	.q_b_18(q_b_181),
	.q_b_17(q_b_171),
	.q_b_31(q_b_312),
	.q_b_30(q_b_301),
	.q_b_29(q_b_291),
	.q_b_28(q_b_281),
	.q_b_27(q_b_271),
	.q_b_26(q_b_261),
	.q_b_25(q_b_251),
	.q_b_10(q_b_101),
	.q_b_24(q_b_241),
	.q_b_9(q_b_91),
	.q_b_23(q_b_231),
	.q_b_8(q_b_81),
	.q_b_22(q_b_221),
	.q_b_7(q_b_71),
	.q_b_6(q_b_61),
	.q_b_20(q_b_201),
	.q_b_19(q_b_191),
	.counter_reg_bit_0(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.full_dff(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.counter_reg_bit_1(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.data_in_shift_reg_0(\data_in_shift_reg[0]~q ),
	.comb(\comb~1_combout ),
	.comb1(\comb~3_combout ),
	.empty_dff(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.comb2(\comb~4_combout ),
	.data_in_shift_reg_1(\data_in_shift_reg[1]~q ),
	.data_in_shift_reg_2(\data_in_shift_reg[2]~q ),
	.data_in_shift_reg_3(\data_in_shift_reg[3]~q ),
	.data_in_shift_reg_4(\data_in_shift_reg[4]~q ),
	.data_in_shift_reg_11(\data_in_shift_reg[11]~q ),
	.data_in_shift_reg_13(\data_in_shift_reg[13]~q ),
	.data_in_shift_reg_16(\data_in_shift_reg[16]~q ),
	.data_in_shift_reg_12(\data_in_shift_reg[12]~q ),
	.data_in_shift_reg_5(\data_in_shift_reg[5]~q ),
	.data_in_shift_reg_14(\data_in_shift_reg[14]~q ),
	.data_in_shift_reg_15(\data_in_shift_reg[15]~q ),
	.data_in_shift_reg_21(\data_in_shift_reg[21]~q ),
	.data_in_shift_reg_18(\data_in_shift_reg[18]~q ),
	.data_in_shift_reg_17(\data_in_shift_reg[17]~q ),
	.data_in_shift_reg_31(\data_in_shift_reg[31]~q ),
	.data_in_shift_reg_30(\data_in_shift_reg[30]~q ),
	.data_in_shift_reg_29(\data_in_shift_reg[29]~q ),
	.data_in_shift_reg_28(\data_in_shift_reg[28]~q ),
	.data_in_shift_reg_27(\data_in_shift_reg[27]~q ),
	.data_in_shift_reg_26(\data_in_shift_reg[26]~q ),
	.data_in_shift_reg_25(\data_in_shift_reg[25]~q ),
	.data_in_shift_reg_10(\data_in_shift_reg[10]~q ),
	.data_in_shift_reg_24(\data_in_shift_reg[24]~q ),
	.data_in_shift_reg_9(\data_in_shift_reg[9]~q ),
	.data_in_shift_reg_23(\data_in_shift_reg[23]~q ),
	.data_in_shift_reg_8(\data_in_shift_reg[8]~q ),
	.data_in_shift_reg_22(\data_in_shift_reg[22]~q ),
	.data_in_shift_reg_7(\data_in_shift_reg[7]~q ),
	.data_in_shift_reg_6(\data_in_shift_reg[6]~q ),
	.data_in_shift_reg_20(\data_in_shift_reg[20]~q ),
	.data_in_shift_reg_19(\data_in_shift_reg[19]~q ),
	.comb3(comb),
	.GND_port(GND_port));

final_project_soc_altera_up_sync_fifo Audio_In_Left_Channel_FIFO(
	.clk_0(clk_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_11(q_b_111),
	.q_b_13(q_b_13),
	.q_b_16(q_b_16),
	.q_b_12(q_b_12),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_21(q_b_211),
	.q_b_18(q_b_18),
	.q_b_17(q_b_17),
	.q_b_31(q_b_311),
	.q_b_30(q_b_30),
	.q_b_29(q_b_29),
	.q_b_28(q_b_28),
	.q_b_27(q_b_27),
	.q_b_26(q_b_26),
	.q_b_25(q_b_25),
	.q_b_10(q_b_10),
	.q_b_24(q_b_24),
	.q_b_9(q_b_9),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_22(q_b_22),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_20(q_b_20),
	.q_b_19(q_b_19),
	.full_dff(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.counter_reg_bit_3(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_5(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_6(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.counter_reg_bit_2(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.comb(\comb~0_combout ),
	.data_in_shift_reg_0(\data_in_shift_reg[0]~q ),
	.comb1(\comb~1_combout ),
	.empty_dff(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.comb2(\comb~2_combout ),
	.data_in_shift_reg_1(\data_in_shift_reg[1]~q ),
	.data_in_shift_reg_2(\data_in_shift_reg[2]~q ),
	.data_in_shift_reg_3(\data_in_shift_reg[3]~q ),
	.data_in_shift_reg_4(\data_in_shift_reg[4]~q ),
	.data_in_shift_reg_11(\data_in_shift_reg[11]~q ),
	.data_in_shift_reg_13(\data_in_shift_reg[13]~q ),
	.data_in_shift_reg_16(\data_in_shift_reg[16]~q ),
	.data_in_shift_reg_12(\data_in_shift_reg[12]~q ),
	.data_in_shift_reg_5(\data_in_shift_reg[5]~q ),
	.data_in_shift_reg_14(\data_in_shift_reg[14]~q ),
	.data_in_shift_reg_15(\data_in_shift_reg[15]~q ),
	.data_in_shift_reg_21(\data_in_shift_reg[21]~q ),
	.data_in_shift_reg_18(\data_in_shift_reg[18]~q ),
	.data_in_shift_reg_17(\data_in_shift_reg[17]~q ),
	.data_in_shift_reg_31(\data_in_shift_reg[31]~q ),
	.data_in_shift_reg_30(\data_in_shift_reg[30]~q ),
	.data_in_shift_reg_29(\data_in_shift_reg[29]~q ),
	.data_in_shift_reg_28(\data_in_shift_reg[28]~q ),
	.data_in_shift_reg_27(\data_in_shift_reg[27]~q ),
	.data_in_shift_reg_26(\data_in_shift_reg[26]~q ),
	.data_in_shift_reg_25(\data_in_shift_reg[25]~q ),
	.data_in_shift_reg_10(\data_in_shift_reg[10]~q ),
	.data_in_shift_reg_24(\data_in_shift_reg[24]~q ),
	.data_in_shift_reg_9(\data_in_shift_reg[9]~q ),
	.data_in_shift_reg_23(\data_in_shift_reg[23]~q ),
	.data_in_shift_reg_8(\data_in_shift_reg[8]~q ),
	.data_in_shift_reg_22(\data_in_shift_reg[22]~q ),
	.data_in_shift_reg_7(\data_in_shift_reg[7]~q ),
	.data_in_shift_reg_6(\data_in_shift_reg[6]~q ),
	.data_in_shift_reg_20(\data_in_shift_reg[20]~q ),
	.data_in_shift_reg_19(\data_in_shift_reg[19]~q ),
	.comb3(comb),
	.GND_port(GND_port));

final_project_soc_altera_up_audio_bit_counter Audio_Out_Bit_Counter(
	.clk(clk_0),
	.counting1(\Audio_Out_Bit_Counter|counting~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.falling_edge(falling_edge),
	.clear_read_fifos(clear_read_fifos),
	.comb(comb),
	.found_edge(found_edge));

cycloneive_lcell_comb \comb~0 (
	.dataa(last_test_clk1),
	.datab(done_adc_channel_sync),
	.datac(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datad(cur_test_clk1),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hEFFF;
defparam \comb~0 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[0] (
	.clk(clk_0),
	.d(\data_in_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[0]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[0] .is_wysiwyg = "true";
defparam \data_in_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \comb~1 (
	.dataa(src_data_39),
	.datab(WideOr1),
	.datac(src_data_68),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'hFDFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~2 (
	.dataa(\comb~1_combout ),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datac(gnd),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
defparam \comb~2 .lut_mask = 16'hEEFF;
defparam \comb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~3 (
	.dataa(cur_test_clk1),
	.datab(done_adc_channel_sync),
	.datac(last_test_clk1),
	.datad(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~3_combout ),
	.cout());
defparam \comb~3 .lut_mask = 16'hEFFF;
defparam \comb~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~4 (
	.dataa(src_data_38),
	.datab(\comb~1_combout ),
	.datac(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\comb~4_combout ),
	.cout());
defparam \comb~4 .lut_mask = 16'hFEFE;
defparam \comb~4 .sum_lutc_input = "datac";

dffeas \data_in_shift_reg[1] (
	.clk(clk_0),
	.d(\data_in_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[1]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[1] .is_wysiwyg = "true";
defparam \data_in_shift_reg[1] .power_up = "low";

dffeas \data_in_shift_reg[2] (
	.clk(clk_0),
	.d(\data_in_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[2]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[2] .is_wysiwyg = "true";
defparam \data_in_shift_reg[2] .power_up = "low";

dffeas \data_in_shift_reg[3] (
	.clk(clk_0),
	.d(\data_in_shift_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[3]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[3] .is_wysiwyg = "true";
defparam \data_in_shift_reg[3] .power_up = "low";

dffeas \data_in_shift_reg[4] (
	.clk(clk_0),
	.d(\data_in_shift_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[4]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[4] .is_wysiwyg = "true";
defparam \data_in_shift_reg[4] .power_up = "low";

dffeas \data_in_shift_reg[11] (
	.clk(clk_0),
	.d(\data_in_shift_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[11]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[11] .is_wysiwyg = "true";
defparam \data_in_shift_reg[11] .power_up = "low";

dffeas \data_in_shift_reg[13] (
	.clk(clk_0),
	.d(\data_in_shift_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[13]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[13] .is_wysiwyg = "true";
defparam \data_in_shift_reg[13] .power_up = "low";

dffeas \data_in_shift_reg[16] (
	.clk(clk_0),
	.d(\data_in_shift_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[16]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[16] .is_wysiwyg = "true";
defparam \data_in_shift_reg[16] .power_up = "low";

dffeas \data_in_shift_reg[12] (
	.clk(clk_0),
	.d(\data_in_shift_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[12]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[12] .is_wysiwyg = "true";
defparam \data_in_shift_reg[12] .power_up = "low";

dffeas \data_in_shift_reg[5] (
	.clk(clk_0),
	.d(\data_in_shift_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[5]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[5] .is_wysiwyg = "true";
defparam \data_in_shift_reg[5] .power_up = "low";

dffeas \data_in_shift_reg[14] (
	.clk(clk_0),
	.d(\data_in_shift_reg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[14]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[14] .is_wysiwyg = "true";
defparam \data_in_shift_reg[14] .power_up = "low";

dffeas \data_in_shift_reg[15] (
	.clk(clk_0),
	.d(\data_in_shift_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[15]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[15] .is_wysiwyg = "true";
defparam \data_in_shift_reg[15] .power_up = "low";

dffeas \data_in_shift_reg[21] (
	.clk(clk_0),
	.d(\data_in_shift_reg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[21]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[21] .is_wysiwyg = "true";
defparam \data_in_shift_reg[21] .power_up = "low";

dffeas \data_in_shift_reg[18] (
	.clk(clk_0),
	.d(\data_in_shift_reg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[18]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[18] .is_wysiwyg = "true";
defparam \data_in_shift_reg[18] .power_up = "low";

dffeas \data_in_shift_reg[17] (
	.clk(clk_0),
	.d(\data_in_shift_reg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[17]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[17] .is_wysiwyg = "true";
defparam \data_in_shift_reg[17] .power_up = "low";

dffeas \data_in_shift_reg[31] (
	.clk(clk_0),
	.d(\data_in_shift_reg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[31]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[31] .is_wysiwyg = "true";
defparam \data_in_shift_reg[31] .power_up = "low";

dffeas \data_in_shift_reg[30] (
	.clk(clk_0),
	.d(\data_in_shift_reg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[30]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[30] .is_wysiwyg = "true";
defparam \data_in_shift_reg[30] .power_up = "low";

dffeas \data_in_shift_reg[29] (
	.clk(clk_0),
	.d(\data_in_shift_reg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[29]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[29] .is_wysiwyg = "true";
defparam \data_in_shift_reg[29] .power_up = "low";

dffeas \data_in_shift_reg[28] (
	.clk(clk_0),
	.d(\data_in_shift_reg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[28]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[28] .is_wysiwyg = "true";
defparam \data_in_shift_reg[28] .power_up = "low";

dffeas \data_in_shift_reg[27] (
	.clk(clk_0),
	.d(\data_in_shift_reg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[27]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[27] .is_wysiwyg = "true";
defparam \data_in_shift_reg[27] .power_up = "low";

dffeas \data_in_shift_reg[26] (
	.clk(clk_0),
	.d(\data_in_shift_reg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[26]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[26] .is_wysiwyg = "true";
defparam \data_in_shift_reg[26] .power_up = "low";

dffeas \data_in_shift_reg[25] (
	.clk(clk_0),
	.d(\data_in_shift_reg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[25]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[25] .is_wysiwyg = "true";
defparam \data_in_shift_reg[25] .power_up = "low";

dffeas \data_in_shift_reg[10] (
	.clk(clk_0),
	.d(\data_in_shift_reg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[10]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[10] .is_wysiwyg = "true";
defparam \data_in_shift_reg[10] .power_up = "low";

dffeas \data_in_shift_reg[24] (
	.clk(clk_0),
	.d(\data_in_shift_reg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[24]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[24] .is_wysiwyg = "true";
defparam \data_in_shift_reg[24] .power_up = "low";

dffeas \data_in_shift_reg[9] (
	.clk(clk_0),
	.d(\data_in_shift_reg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[9]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[9] .is_wysiwyg = "true";
defparam \data_in_shift_reg[9] .power_up = "low";

dffeas \data_in_shift_reg[23] (
	.clk(clk_0),
	.d(\data_in_shift_reg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[23]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[23] .is_wysiwyg = "true";
defparam \data_in_shift_reg[23] .power_up = "low";

dffeas \data_in_shift_reg[8] (
	.clk(clk_0),
	.d(\data_in_shift_reg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[8]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[8] .is_wysiwyg = "true";
defparam \data_in_shift_reg[8] .power_up = "low";

dffeas \data_in_shift_reg[22] (
	.clk(clk_0),
	.d(\data_in_shift_reg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[22]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[22] .is_wysiwyg = "true";
defparam \data_in_shift_reg[22] .power_up = "low";

dffeas \data_in_shift_reg[7] (
	.clk(clk_0),
	.d(\data_in_shift_reg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[7]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[7] .is_wysiwyg = "true";
defparam \data_in_shift_reg[7] .power_up = "low";

dffeas \data_in_shift_reg[6] (
	.clk(clk_0),
	.d(\data_in_shift_reg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[6]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[6] .is_wysiwyg = "true";
defparam \data_in_shift_reg[6] .power_up = "low";

dffeas \data_in_shift_reg[20] (
	.clk(clk_0),
	.d(\data_in_shift_reg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[20]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[20] .is_wysiwyg = "true";
defparam \data_in_shift_reg[20] .power_up = "low";

dffeas \data_in_shift_reg[19] (
	.clk(clk_0),
	.d(\data_in_shift_reg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_in_shift_reg[9]~1_combout ),
	.q(\data_in_shift_reg[19]~q ),
	.prn(vcc));
defparam \data_in_shift_reg[19] .is_wysiwyg = "true";
defparam \data_in_shift_reg[19] .power_up = "low";

cycloneive_lcell_comb \data_in_shift_reg~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(audio_wire_ADCDAT),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~0_combout ),
	.cout());
defparam \data_in_shift_reg~0 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg[9]~1 (
	.dataa(comb),
	.datab(last_test_clk),
	.datac(cur_test_clk),
	.datad(\Audio_Out_Bit_Counter|counting~q ),
	.cin(gnd),
	.combout(\data_in_shift_reg[9]~1_combout ),
	.cout());
defparam \data_in_shift_reg[9]~1 .lut_mask = 16'hFFFB;
defparam \data_in_shift_reg[9]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[0]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~2_combout ),
	.cout());
defparam \data_in_shift_reg~2 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[1]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~3_combout ),
	.cout());
defparam \data_in_shift_reg~3 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[2]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~4_combout ),
	.cout());
defparam \data_in_shift_reg~4 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[3]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~5_combout ),
	.cout());
defparam \data_in_shift_reg~5 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[10]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~6_combout ),
	.cout());
defparam \data_in_shift_reg~6 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[12]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~7_combout ),
	.cout());
defparam \data_in_shift_reg~7 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~8 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[15]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~8_combout ),
	.cout());
defparam \data_in_shift_reg~8 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~9 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[11]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~9_combout ),
	.cout());
defparam \data_in_shift_reg~9 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~10 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[4]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~10_combout ),
	.cout());
defparam \data_in_shift_reg~10 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~11 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[13]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~11_combout ),
	.cout());
defparam \data_in_shift_reg~11 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~12 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[14]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~12_combout ),
	.cout());
defparam \data_in_shift_reg~12 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~13 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[20]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~13_combout ),
	.cout());
defparam \data_in_shift_reg~13 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~14 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[17]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~14_combout ),
	.cout());
defparam \data_in_shift_reg~14 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~15 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[16]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~15_combout ),
	.cout());
defparam \data_in_shift_reg~15 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~16 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[30]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~16_combout ),
	.cout());
defparam \data_in_shift_reg~16 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~17 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[29]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~17_combout ),
	.cout());
defparam \data_in_shift_reg~17 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~18 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[28]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~18_combout ),
	.cout());
defparam \data_in_shift_reg~18 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~19 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[27]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~19_combout ),
	.cout());
defparam \data_in_shift_reg~19 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~20 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[26]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~20_combout ),
	.cout());
defparam \data_in_shift_reg~20 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~21 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[25]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~21_combout ),
	.cout());
defparam \data_in_shift_reg~21 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~22 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[24]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~22_combout ),
	.cout());
defparam \data_in_shift_reg~22 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~23 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[9]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~23_combout ),
	.cout());
defparam \data_in_shift_reg~23 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~24 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[23]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~24_combout ),
	.cout());
defparam \data_in_shift_reg~24 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~25 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[8]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~25_combout ),
	.cout());
defparam \data_in_shift_reg~25 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~26 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[22]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~26_combout ),
	.cout());
defparam \data_in_shift_reg~26 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~27 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[7]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~27_combout ),
	.cout());
defparam \data_in_shift_reg~27 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~28 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[21]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~28_combout ),
	.cout());
defparam \data_in_shift_reg~28 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~29 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[6]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~29_combout ),
	.cout());
defparam \data_in_shift_reg~29 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[5]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~30_combout ),
	.cout());
defparam \data_in_shift_reg~30 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[19]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~31_combout ),
	.cout());
defparam \data_in_shift_reg~31 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_shift_reg~32 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\data_in_shift_reg[18]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\data_in_shift_reg~32_combout ),
	.cout());
defparam \data_in_shift_reg~32 .lut_mask = 16'hEEFF;
defparam \data_in_shift_reg~32 .sum_lutc_input = "datac";

dffeas \right_audio_fifo_read_space[0] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_0),
	.prn(vcc));
defparam \right_audio_fifo_read_space[0] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[0] .power_up = "low";

dffeas \right_audio_fifo_read_space[1] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_1),
	.prn(vcc));
defparam \right_audio_fifo_read_space[1] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[1] .power_up = "low";

dffeas \right_audio_fifo_read_space[2] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_2),
	.prn(vcc));
defparam \right_audio_fifo_read_space[2] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[2] .power_up = "low";

dffeas \right_audio_fifo_read_space[3] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_3),
	.prn(vcc));
defparam \right_audio_fifo_read_space[3] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[3] .power_up = "low";

dffeas \right_audio_fifo_read_space[4] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_4),
	.prn(vcc));
defparam \right_audio_fifo_read_space[4] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[4] .power_up = "low";

dffeas \left_audio_fifo_read_space[3] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_3),
	.prn(vcc));
defparam \left_audio_fifo_read_space[3] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[3] .power_up = "low";

dffeas \left_audio_fifo_read_space[5] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_5),
	.prn(vcc));
defparam \left_audio_fifo_read_space[5] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[5] .power_up = "low";

dffeas \left_audio_fifo_read_space[4] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_4),
	.prn(vcc));
defparam \left_audio_fifo_read_space[4] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[4] .power_up = "low";

dffeas \right_audio_fifo_read_space[5] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_5),
	.prn(vcc));
defparam \right_audio_fifo_read_space[5] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[5] .power_up = "low";

dffeas \left_audio_fifo_read_space[6] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_6),
	.prn(vcc));
defparam \left_audio_fifo_read_space[6] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[6] .power_up = "low";

dffeas \left_audio_fifo_read_space[7] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_7),
	.prn(vcc));
defparam \left_audio_fifo_read_space[7] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[7] .power_up = "low";

dffeas \left_audio_fifo_read_space[2] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_2),
	.prn(vcc));
defparam \left_audio_fifo_read_space[2] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[2] .power_up = "low";

dffeas \left_audio_fifo_read_space[1] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_1),
	.prn(vcc));
defparam \left_audio_fifo_read_space[1] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[1] .power_up = "low";

dffeas \left_audio_fifo_read_space[0] (
	.clk(clk_0),
	.d(\left_audio_fifo_read_space~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(left_audio_fifo_read_space_0),
	.prn(vcc));
defparam \left_audio_fifo_read_space[0] .is_wysiwyg = "true";
defparam \left_audio_fifo_read_space[0] .power_up = "low";

dffeas \right_audio_fifo_read_space[7] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_7),
	.prn(vcc));
defparam \right_audio_fifo_read_space[7] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[7] .power_up = "low";

dffeas \right_audio_fifo_read_space[6] (
	.clk(clk_0),
	.d(\right_audio_fifo_read_space~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(right_audio_fifo_read_space_6),
	.prn(vcc));
defparam \right_audio_fifo_read_space[6] .is_wysiwyg = "true";
defparam \right_audio_fifo_read_space[6] .power_up = "low";

cycloneive_lcell_comb \right_audio_fifo_read_space~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~0_combout ),
	.cout());
defparam \right_audio_fifo_read_space~0 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~1_combout ),
	.cout());
defparam \right_audio_fifo_read_space~1 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~2_combout ),
	.cout());
defparam \right_audio_fifo_read_space~2 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~3_combout ),
	.cout());
defparam \right_audio_fifo_read_space~3 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~4_combout ),
	.cout());
defparam \right_audio_fifo_read_space~4 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~0_combout ),
	.cout());
defparam \left_audio_fifo_read_space~0 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~1 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~1_combout ),
	.cout());
defparam \left_audio_fifo_read_space~1 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~2_combout ),
	.cout());
defparam \left_audio_fifo_read_space~2 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~5_combout ),
	.cout());
defparam \right_audio_fifo_read_space~5 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~3_combout ),
	.cout());
defparam \left_audio_fifo_read_space~3 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~4_combout ),
	.cout());
defparam \left_audio_fifo_read_space~4 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~5_combout ),
	.cout());
defparam \left_audio_fifo_read_space~5 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~6_combout ),
	.cout());
defparam \left_audio_fifo_read_space~6 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_audio_fifo_read_space~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\left_audio_fifo_read_space~7_combout ),
	.cout());
defparam \left_audio_fifo_read_space~7 .lut_mask = 16'hEEFF;
defparam \left_audio_fifo_read_space~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~6 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~6_combout ),
	.cout());
defparam \right_audio_fifo_read_space~6 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_audio_fifo_read_space~7 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\Audio_In_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datac(gnd),
	.datad(clear_read_fifos),
	.cin(gnd),
	.combout(\right_audio_fifo_read_space~7_combout ),
	.cout());
defparam \right_audio_fifo_read_space~7 .lut_mask = 16'hEEFF;
defparam \right_audio_fifo_read_space~7 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_audio_bit_counter (
	clk,
	counting1,
	altera_reset_synchronizer_int_chain_out,
	falling_edge,
	clear_read_fifos,
	comb,
	found_edge)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	counting1;
input 	altera_reset_synchronizer_int_chain_out;
input 	falling_edge;
input 	clear_read_fifos;
input 	comb;
input 	found_edge;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~20_combout ;
wire \Add0~30_combout ;
wire \bit_counter[3]~2_combout ;
wire \bit_counter[0]~q ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \Add0~31_combout ;
wire \bit_counter[1]~q ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \Add0~32_combout ;
wire \bit_counter[2]~q ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \Add0~33_combout ;
wire \bit_counter[3]~q ;
wire \bit_counter[3]~0_combout ;
wire \Add0~27 ;
wire \Add0~28_combout ;
wire \Add0~34_combout ;
wire \bit_counter[4]~q ;
wire \bit_counter[3]~1_combout ;
wire \counting~0_combout ;


dffeas counting(
	.clk(clk),
	.d(\counting~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(counting1),
	.prn(vcc));
defparam counting.is_wysiwyg = "true";
defparam counting.power_up = "low";

cycloneive_lcell_comb \Add0~20 (
	.dataa(\bit_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h55AA;
defparam \Add0~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~30 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(found_edge),
	.datad(\Add0~20_combout ),
	.cin(gnd),
	.combout(\Add0~30_combout ),
	.cout());
defparam \Add0~30 .lut_mask = 16'hFFFB;
defparam \Add0~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \bit_counter[3]~2 (
	.dataa(comb),
	.datab(falling_edge),
	.datac(\bit_counter[3]~1_combout ),
	.datad(found_edge),
	.cin(gnd),
	.combout(\bit_counter[3]~2_combout ),
	.cout());
defparam \bit_counter[3]~2 .lut_mask = 16'hFFBF;
defparam \bit_counter[3]~2 .sum_lutc_input = "datac";

dffeas \bit_counter[0] (
	.clk(clk),
	.d(\Add0~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bit_counter[3]~2_combout ),
	.q(\bit_counter[0]~q ),
	.prn(vcc));
defparam \bit_counter[0] .is_wysiwyg = "true";
defparam \bit_counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~22 (
	.dataa(\bit_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~31 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(found_edge),
	.datad(\Add0~22_combout ),
	.cin(gnd),
	.combout(\Add0~31_combout ),
	.cout());
defparam \Add0~31 .lut_mask = 16'hFFFB;
defparam \Add0~31 .sum_lutc_input = "datac";

dffeas \bit_counter[1] (
	.clk(clk),
	.d(\Add0~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bit_counter[3]~2_combout ),
	.q(\bit_counter[1]~q ),
	.prn(vcc));
defparam \bit_counter[1] .is_wysiwyg = "true";
defparam \bit_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add0~24 (
	.dataa(\bit_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'h5AAF;
defparam \Add0~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~32 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(found_edge),
	.datad(\Add0~24_combout ),
	.cin(gnd),
	.combout(\Add0~32_combout ),
	.cout());
defparam \Add0~32 .lut_mask = 16'hFFFB;
defparam \Add0~32 .sum_lutc_input = "datac";

dffeas \bit_counter[2] (
	.clk(clk),
	.d(\Add0~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bit_counter[3]~2_combout ),
	.q(\bit_counter[2]~q ),
	.prn(vcc));
defparam \bit_counter[2] .is_wysiwyg = "true";
defparam \bit_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add0~26 (
	.dataa(\bit_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
defparam \Add0~26 .lut_mask = 16'h5A5F;
defparam \Add0~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~33 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(found_edge),
	.datad(\Add0~26_combout ),
	.cin(gnd),
	.combout(\Add0~33_combout ),
	.cout());
defparam \Add0~33 .lut_mask = 16'hFFFB;
defparam \Add0~33 .sum_lutc_input = "datac";

dffeas \bit_counter[3] (
	.clk(clk),
	.d(\Add0~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bit_counter[3]~2_combout ),
	.q(\bit_counter[3]~q ),
	.prn(vcc));
defparam \bit_counter[3] .is_wysiwyg = "true";
defparam \bit_counter[3] .power_up = "low";

cycloneive_lcell_comb \bit_counter[3]~0 (
	.dataa(\bit_counter[0]~q ),
	.datab(\bit_counter[1]~q ),
	.datac(\bit_counter[2]~q ),
	.datad(\bit_counter[3]~q ),
	.cin(gnd),
	.combout(\bit_counter[3]~0_combout ),
	.cout());
defparam \bit_counter[3]~0 .lut_mask = 16'h7FFF;
defparam \bit_counter[3]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~28 (
	.dataa(\bit_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout());
defparam \Add0~28 .lut_mask = 16'h5A5A;
defparam \Add0~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~34 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(found_edge),
	.datad(\Add0~28_combout ),
	.cin(gnd),
	.combout(\Add0~34_combout ),
	.cout());
defparam \Add0~34 .lut_mask = 16'hFFFB;
defparam \Add0~34 .sum_lutc_input = "datac";

dffeas \bit_counter[4] (
	.clk(clk),
	.d(\Add0~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bit_counter[3]~2_combout ),
	.q(\bit_counter[4]~q ),
	.prn(vcc));
defparam \bit_counter[4] .is_wysiwyg = "true";
defparam \bit_counter[4] .power_up = "low";

cycloneive_lcell_comb \bit_counter[3]~1 (
	.dataa(\bit_counter[3]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\bit_counter[4]~q ),
	.cin(gnd),
	.combout(\bit_counter[3]~1_combout ),
	.cout());
defparam \bit_counter[3]~1 .lut_mask = 16'hAAFF;
defparam \bit_counter[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counting~0 (
	.dataa(found_edge),
	.datab(counting1),
	.datac(falling_edge),
	.datad(\bit_counter[3]~1_combout ),
	.cin(gnd),
	.combout(\counting~0_combout ),
	.cout());
defparam \counting~0 .lut_mask = 16'hFEFF;
defparam \counting~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_sync_fifo (
	clk_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_11,
	q_b_13,
	q_b_16,
	q_b_12,
	q_b_5,
	q_b_14,
	q_b_15,
	q_b_21,
	q_b_18,
	q_b_17,
	q_b_31,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_10,
	q_b_24,
	q_b_9,
	q_b_23,
	q_b_8,
	q_b_22,
	q_b_7,
	q_b_6,
	q_b_20,
	q_b_19,
	full_dff,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	comb,
	data_in_shift_reg_0,
	comb1,
	empty_dff,
	comb2,
	data_in_shift_reg_1,
	data_in_shift_reg_2,
	data_in_shift_reg_3,
	data_in_shift_reg_4,
	data_in_shift_reg_11,
	data_in_shift_reg_13,
	data_in_shift_reg_16,
	data_in_shift_reg_12,
	data_in_shift_reg_5,
	data_in_shift_reg_14,
	data_in_shift_reg_15,
	data_in_shift_reg_21,
	data_in_shift_reg_18,
	data_in_shift_reg_17,
	data_in_shift_reg_31,
	data_in_shift_reg_30,
	data_in_shift_reg_29,
	data_in_shift_reg_28,
	data_in_shift_reg_27,
	data_in_shift_reg_26,
	data_in_shift_reg_25,
	data_in_shift_reg_10,
	data_in_shift_reg_24,
	data_in_shift_reg_9,
	data_in_shift_reg_23,
	data_in_shift_reg_8,
	data_in_shift_reg_22,
	data_in_shift_reg_7,
	data_in_shift_reg_6,
	data_in_shift_reg_20,
	data_in_shift_reg_19,
	comb3,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_11;
output 	q_b_13;
output 	q_b_16;
output 	q_b_12;
output 	q_b_5;
output 	q_b_14;
output 	q_b_15;
output 	q_b_21;
output 	q_b_18;
output 	q_b_17;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_10;
output 	q_b_24;
output 	q_b_9;
output 	q_b_23;
output 	q_b_8;
output 	q_b_22;
output 	q_b_7;
output 	q_b_6;
output 	q_b_20;
output 	q_b_19;
output 	full_dff;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	comb;
input 	data_in_shift_reg_0;
input 	comb1;
output 	empty_dff;
input 	comb2;
input 	data_in_shift_reg_1;
input 	data_in_shift_reg_2;
input 	data_in_shift_reg_3;
input 	data_in_shift_reg_4;
input 	data_in_shift_reg_11;
input 	data_in_shift_reg_13;
input 	data_in_shift_reg_16;
input 	data_in_shift_reg_12;
input 	data_in_shift_reg_5;
input 	data_in_shift_reg_14;
input 	data_in_shift_reg_15;
input 	data_in_shift_reg_21;
input 	data_in_shift_reg_18;
input 	data_in_shift_reg_17;
input 	data_in_shift_reg_31;
input 	data_in_shift_reg_30;
input 	data_in_shift_reg_29;
input 	data_in_shift_reg_28;
input 	data_in_shift_reg_27;
input 	data_in_shift_reg_26;
input 	data_in_shift_reg_25;
input 	data_in_shift_reg_10;
input 	data_in_shift_reg_24;
input 	data_in_shift_reg_9;
input 	data_in_shift_reg_23;
input 	data_in_shift_reg_8;
input 	data_in_shift_reg_22;
input 	data_in_shift_reg_7;
input 	data_in_shift_reg_6;
input 	data_in_shift_reg_20;
input 	data_in_shift_reg_19;
input 	comb3;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_1 Sync_FIFO(
	.clock(clk_0),
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.full_dff(full_dff),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.wrreq(comb),
	.data({data_in_shift_reg_31,data_in_shift_reg_30,data_in_shift_reg_29,data_in_shift_reg_28,data_in_shift_reg_27,data_in_shift_reg_26,data_in_shift_reg_25,data_in_shift_reg_24,data_in_shift_reg_23,data_in_shift_reg_22,data_in_shift_reg_21,data_in_shift_reg_20,
data_in_shift_reg_19,data_in_shift_reg_18,data_in_shift_reg_17,data_in_shift_reg_16,data_in_shift_reg_15,data_in_shift_reg_14,data_in_shift_reg_13,data_in_shift_reg_12,data_in_shift_reg_11,data_in_shift_reg_10,data_in_shift_reg_9,data_in_shift_reg_8,
data_in_shift_reg_7,data_in_shift_reg_6,data_in_shift_reg_5,data_in_shift_reg_4,data_in_shift_reg_3,data_in_shift_reg_2,data_in_shift_reg_1,data_in_shift_reg_0}),
	.comb(comb1),
	.empty_dff(empty_dff),
	.comb1(comb2),
	.comb2(comb3),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_1 (
	clock,
	q,
	full_dff,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	wrreq,
	data,
	comb,
	empty_dff,
	comb1,
	comb2,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	full_dff;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	wrreq;
input 	[31:0] data;
input 	comb;
output 	empty_dff;
input 	comb1;
input 	comb2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_n441 auto_generated(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.full_dff(full_dff),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.wrreq(wrreq),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.empty_dff(empty_dff),
	.comb1(comb1),
	.comb2(comb2),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_n441 (
	clock,
	q,
	full_dff,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	wrreq,
	data,
	comb,
	empty_dff,
	comb1,
	comb2,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	full_dff;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	wrreq;
input 	[31:0] data;
input 	comb;
output 	empty_dff;
input 	comb1;
input 	comb2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_a_dpfifo_as31 dpfifo(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.full_dff1(full_dff),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.wreq(wrreq),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.empty_dff1(empty_dff),
	.comb1(comb1),
	.comb2(comb2),
	.GND_port(GND_port));

endmodule

module final_project_soc_a_dpfifo_as31 (
	clock,
	q,
	full_dff1,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	wreq,
	data,
	comb,
	empty_dff1,
	comb1,
	comb2,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	full_dff1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	wreq;
input 	[31:0] data;
input 	comb;
output 	empty_dff1;
input 	comb1;
input 	comb2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_2~0_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_0~2_combout ;
wire \usedw_will_be_0~3_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~3_combout ;
wire \usedw_will_be_1~4_combout ;
wire \empty_dff~0_combout ;


final_project_soc_cntr_0ab wr_ptr(
	.clock(clock),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_read_fifos(clear_read_fifos),
	.comb(wreq),
	.comb1(comb2),
	.GND_port(GND_port));

final_project_soc_cntr_ca7 usedw_counter(
	.clock(clock),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_read_fifos(clear_read_fifos),
	.updown(wreq),
	.comb(comb1),
	.comb1(comb2),
	.GND_port(GND_port));

final_project_soc_cntr_v9b rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_read_fifos(clear_read_fifos),
	.comb(comb1),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.comb1(comb2),
	.GND_port(GND_port));

final_project_soc_altsyncram_dh81 FIFOram(
	.clock0(clock),
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(wreq),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(comb1),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(comb2),
	.datab(\low_addressa[0]~q ),
	.datac(comb1),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hC5FF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(clear_read_fifos),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hFF77;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(comb),
	.datab(empty_dff1),
	.datac(src_data_38),
	.datad(comb2),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hFFEF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hDDF5;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hDDF5;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hDDF5;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hDDF5;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datac(\low_addressa[5]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hDDF5;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datac(\low_addressa[6]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hDDF5;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb2),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_6),
	.datac(counter_reg_bit_0),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_3),
	.datac(counter_reg_bit_4),
	.datad(\_~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(full_dff1),
	.datab(wreq),
	.datac(\_~1_combout ),
	.datad(comb1),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_6),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hEFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(\_~3_combout ),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hBFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~0_combout ),
	.datab(comb1),
	.datac(\_~4_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb2),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(comb1),
	.datab(\usedw_is_2_dff~q ),
	.datac(gnd),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hEEFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~2 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\usedw_will_be_0~2_combout ),
	.cout());
defparam \usedw_will_be_0~2 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(\usedw_will_be_0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_0~3_combout ),
	.cout());
defparam \usedw_will_be_0~3 .lut_mask = 16'hFBFB;
defparam \usedw_will_be_0~3 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(comb1),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hFFFB;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(wreq),
	.datab(\usedw_will_be_1~4_combout ),
	.datac(comb2),
	.datad(\usedw_will_be_0~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altsyncram_dh81 (
	clock0,
	q_b,
	address_a,
	wren_a,
	data_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[6:0] address_a;
input 	wren_a;
input 	[31:0] data_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 7;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 127;
defparam ram_block1a16.port_a_logical_ram_depth = 128;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 7;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 127;
defparam ram_block1a16.port_b_logical_ram_depth = 128;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 7;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 127;
defparam ram_block1a21.port_a_logical_ram_depth = 128;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 7;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 127;
defparam ram_block1a21.port_b_logical_ram_depth = 128;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 7;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 127;
defparam ram_block1a18.port_a_logical_ram_depth = 128;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 7;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 127;
defparam ram_block1a18.port_b_logical_ram_depth = 128;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 7;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 127;
defparam ram_block1a17.port_a_logical_ram_depth = 128;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 7;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 127;
defparam ram_block1a17.port_b_logical_ram_depth = 128;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 7;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 127;
defparam ram_block1a31.port_a_logical_ram_depth = 128;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 7;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 127;
defparam ram_block1a31.port_b_logical_ram_depth = 128;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 7;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 127;
defparam ram_block1a30.port_a_logical_ram_depth = 128;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 7;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 127;
defparam ram_block1a30.port_b_logical_ram_depth = 128;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 7;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 127;
defparam ram_block1a29.port_a_logical_ram_depth = 128;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 7;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 127;
defparam ram_block1a29.port_b_logical_ram_depth = 128;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 7;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 127;
defparam ram_block1a28.port_a_logical_ram_depth = 128;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 7;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 127;
defparam ram_block1a28.port_b_logical_ram_depth = 128;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 7;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 127;
defparam ram_block1a27.port_a_logical_ram_depth = 128;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 7;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 127;
defparam ram_block1a27.port_b_logical_ram_depth = 128;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 7;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 127;
defparam ram_block1a26.port_a_logical_ram_depth = 128;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 7;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 127;
defparam ram_block1a26.port_b_logical_ram_depth = 128;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 7;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 127;
defparam ram_block1a25.port_a_logical_ram_depth = 128;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 7;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 127;
defparam ram_block1a25.port_b_logical_ram_depth = 128;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 7;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 127;
defparam ram_block1a24.port_a_logical_ram_depth = 128;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 7;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 127;
defparam ram_block1a24.port_b_logical_ram_depth = 128;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 7;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 127;
defparam ram_block1a23.port_a_logical_ram_depth = 128;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 7;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 127;
defparam ram_block1a23.port_b_logical_ram_depth = 128;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 7;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 127;
defparam ram_block1a22.port_a_logical_ram_depth = 128;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 7;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 127;
defparam ram_block1a22.port_b_logical_ram_depth = 128;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 7;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 127;
defparam ram_block1a20.port_a_logical_ram_depth = 128;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 7;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 127;
defparam ram_block1a20.port_b_logical_ram_depth = 128;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 7;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 127;
defparam ram_block1a19.port_a_logical_ram_depth = 128;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 7;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 127;
defparam ram_block1a19.port_b_logical_ram_depth = 128;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

endmodule

module final_project_soc_cntr_0ab (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	clear_read_fifos,
	comb,
	comb1,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_read_fifos;
input 	comb;
input 	comb1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(comb),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFDFD;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_ca7 (
	clock,
	counter_reg_bit_3,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_6,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	altera_reset_synchronizer_int_chain_out,
	clear_read_fifos,
	updown,
	comb,
	comb1,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_3;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_6;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_read_fifos;
input 	updown;
input 	comb;
input 	comb1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \_~2_combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(updown),
	.datad(comb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hDFFD;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_v9b (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	altera_reset_synchronizer_int_chain_out,
	clear_read_fifos,
	comb,
	rd_ptr_lsb,
	comb1,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_read_fifos;
input 	comb;
input 	rd_ptr_lsb;
input 	comb1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(comb),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFDFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_altera_up_sync_fifo_1 (
	clk_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_11,
	q_b_13,
	q_b_16,
	q_b_12,
	q_b_5,
	q_b_14,
	q_b_15,
	q_b_21,
	q_b_18,
	q_b_17,
	q_b_31,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_10,
	q_b_24,
	q_b_9,
	q_b_23,
	q_b_8,
	q_b_22,
	q_b_7,
	q_b_6,
	q_b_20,
	q_b_19,
	counter_reg_bit_0,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	data_in_shift_reg_0,
	comb,
	comb1,
	empty_dff,
	comb2,
	data_in_shift_reg_1,
	data_in_shift_reg_2,
	data_in_shift_reg_3,
	data_in_shift_reg_4,
	data_in_shift_reg_11,
	data_in_shift_reg_13,
	data_in_shift_reg_16,
	data_in_shift_reg_12,
	data_in_shift_reg_5,
	data_in_shift_reg_14,
	data_in_shift_reg_15,
	data_in_shift_reg_21,
	data_in_shift_reg_18,
	data_in_shift_reg_17,
	data_in_shift_reg_31,
	data_in_shift_reg_30,
	data_in_shift_reg_29,
	data_in_shift_reg_28,
	data_in_shift_reg_27,
	data_in_shift_reg_26,
	data_in_shift_reg_25,
	data_in_shift_reg_10,
	data_in_shift_reg_24,
	data_in_shift_reg_9,
	data_in_shift_reg_23,
	data_in_shift_reg_8,
	data_in_shift_reg_22,
	data_in_shift_reg_7,
	data_in_shift_reg_6,
	data_in_shift_reg_20,
	data_in_shift_reg_19,
	comb3,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_11;
output 	q_b_13;
output 	q_b_16;
output 	q_b_12;
output 	q_b_5;
output 	q_b_14;
output 	q_b_15;
output 	q_b_21;
output 	q_b_18;
output 	q_b_17;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_10;
output 	q_b_24;
output 	q_b_9;
output 	q_b_23;
output 	q_b_8;
output 	q_b_22;
output 	q_b_7;
output 	q_b_6;
output 	q_b_20;
output 	q_b_19;
output 	counter_reg_bit_0;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	data_in_shift_reg_0;
input 	comb;
input 	comb1;
output 	empty_dff;
input 	comb2;
input 	data_in_shift_reg_1;
input 	data_in_shift_reg_2;
input 	data_in_shift_reg_3;
input 	data_in_shift_reg_4;
input 	data_in_shift_reg_11;
input 	data_in_shift_reg_13;
input 	data_in_shift_reg_16;
input 	data_in_shift_reg_12;
input 	data_in_shift_reg_5;
input 	data_in_shift_reg_14;
input 	data_in_shift_reg_15;
input 	data_in_shift_reg_21;
input 	data_in_shift_reg_18;
input 	data_in_shift_reg_17;
input 	data_in_shift_reg_31;
input 	data_in_shift_reg_30;
input 	data_in_shift_reg_29;
input 	data_in_shift_reg_28;
input 	data_in_shift_reg_27;
input 	data_in_shift_reg_26;
input 	data_in_shift_reg_25;
input 	data_in_shift_reg_10;
input 	data_in_shift_reg_24;
input 	data_in_shift_reg_9;
input 	data_in_shift_reg_23;
input 	data_in_shift_reg_8;
input 	data_in_shift_reg_22;
input 	data_in_shift_reg_7;
input 	data_in_shift_reg_6;
input 	data_in_shift_reg_20;
input 	data_in_shift_reg_19;
input 	comb3;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_2 Sync_FIFO(
	.clock(clk_0),
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.counter_reg_bit_0(counter_reg_bit_0),
	.full_dff(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_6(counter_reg_bit_6),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.data({data_in_shift_reg_31,data_in_shift_reg_30,data_in_shift_reg_29,data_in_shift_reg_28,data_in_shift_reg_27,data_in_shift_reg_26,data_in_shift_reg_25,data_in_shift_reg_24,data_in_shift_reg_23,data_in_shift_reg_22,data_in_shift_reg_21,data_in_shift_reg_20,
data_in_shift_reg_19,data_in_shift_reg_18,data_in_shift_reg_17,data_in_shift_reg_16,data_in_shift_reg_15,data_in_shift_reg_14,data_in_shift_reg_13,data_in_shift_reg_12,data_in_shift_reg_11,data_in_shift_reg_10,data_in_shift_reg_9,data_in_shift_reg_8,
data_in_shift_reg_7,data_in_shift_reg_6,data_in_shift_reg_5,data_in_shift_reg_4,data_in_shift_reg_3,data_in_shift_reg_2,data_in_shift_reg_1,data_in_shift_reg_0}),
	.comb(comb),
	.wrreq(comb1),
	.empty_dff(empty_dff),
	.comb1(comb2),
	.comb2(comb3),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_2 (
	clock,
	q,
	counter_reg_bit_0,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	data,
	comb,
	wrreq,
	empty_dff,
	comb1,
	comb2,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_0;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	[31:0] data;
input 	comb;
input 	wrreq;
output 	empty_dff;
input 	comb1;
input 	comb2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_n441_1 auto_generated(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_0(counter_reg_bit_0),
	.full_dff(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_6(counter_reg_bit_6),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.wrreq(wrreq),
	.empty_dff(empty_dff),
	.comb1(comb1),
	.comb2(comb2),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_n441_1 (
	clock,
	q,
	counter_reg_bit_0,
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	data,
	comb,
	wrreq,
	empty_dff,
	comb1,
	comb2,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_0;
output 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	[31:0] data;
input 	comb;
input 	wrreq;
output 	empty_dff;
input 	comb1;
input 	comb2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_a_dpfifo_as31_1 dpfifo(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_0(counter_reg_bit_0),
	.full_dff1(full_dff),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_6(counter_reg_bit_6),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_data_38(src_data_38),
	.clear_read_fifos(clear_read_fifos),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.comb(comb),
	.wreq(wrreq),
	.empty_dff1(empty_dff),
	.comb1(comb1),
	.comb2(comb2),
	.GND_port(GND_port));

endmodule

module final_project_soc_a_dpfifo_as31_1 (
	clock,
	q,
	counter_reg_bit_0,
	full_dff1,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	src_data_38,
	clear_read_fifos,
	data,
	comb,
	wreq,
	empty_dff1,
	comb1,
	comb2,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_0;
output 	full_dff1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_data_38;
input 	clear_read_fifos;
input 	[31:0] data;
input 	comb;
input 	wreq;
output 	empty_dff1;
input 	comb1;
input 	comb2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_2~0_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_0~2_combout ;
wire \usedw_will_be_0~3_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~3_combout ;
wire \usedw_will_be_1~4_combout ;
wire \empty_dff~0_combout ;


final_project_soc_cntr_0ab_1 wr_ptr(
	.clock(clock),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_read_fifos(clear_read_fifos),
	.comb(wreq),
	.comb1(comb2),
	.GND_port(GND_port));

final_project_soc_cntr_ca7_1 usedw_counter(
	.clock(clock),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_6(counter_reg_bit_6),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_read_fifos(clear_read_fifos),
	.updown(wreq),
	.comb(comb1),
	.comb1(comb2),
	.GND_port(GND_port));

final_project_soc_cntr_v9b_1 rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_read_fifos(clear_read_fifos),
	.comb(comb1),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.comb1(comb2),
	.GND_port(GND_port));

final_project_soc_altsyncram_dh81_1 FIFOram(
	.clock0(clock),
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(comb1),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(comb2),
	.datab(\low_addressa[0]~q ),
	.datac(comb1),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hC5FF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(clear_read_fifos),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hFF77;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(src_data_38),
	.datab(comb),
	.datac(empty_dff1),
	.datad(comb2),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hFFFE;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hDDF5;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hDDF5;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hDDF5;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hDDF5;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datac(\low_addressa[5]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hDDF5;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(comb2),
	.datab(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datac(\low_addressa[6]~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hDDF5;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb2),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_6),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(counter_reg_bit_4),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_3),
	.datad(\_~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(full_dff1),
	.datab(wreq),
	.datac(\_~1_combout ),
	.datad(comb1),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_6),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hEFFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(\_~3_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hBFFF;
defparam \_~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~0_combout ),
	.datab(comb1),
	.datac(\_~4_combout ),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb2),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(comb1),
	.datab(\usedw_is_2_dff~q ),
	.datac(gnd),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hEEFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~2 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(comb1),
	.cin(gnd),
	.combout(\usedw_will_be_0~2_combout ),
	.cout());
defparam \usedw_will_be_0~2 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(\usedw_will_be_0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_0~3_combout ),
	.cout());
defparam \usedw_will_be_0~3 .lut_mask = 16'hFBFB;
defparam \usedw_will_be_0~3 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(comb1),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~4 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~4_combout ),
	.cout());
defparam \usedw_will_be_1~4 .lut_mask = 16'hFFFB;
defparam \usedw_will_be_1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(wreq),
	.datab(\usedw_will_be_1~4_combout ),
	.datac(comb2),
	.datad(\usedw_will_be_0~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altsyncram_dh81_1 (
	clock0,
	q_b,
	address_a,
	data_a,
	wren_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[6:0] address_a;
input 	[31:0] data_a;
input 	wren_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 7;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 127;
defparam ram_block1a16.port_a_logical_ram_depth = 128;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 7;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 127;
defparam ram_block1a16.port_b_logical_ram_depth = 128;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 7;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 127;
defparam ram_block1a21.port_a_logical_ram_depth = 128;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 7;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 127;
defparam ram_block1a21.port_b_logical_ram_depth = 128;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 7;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 127;
defparam ram_block1a18.port_a_logical_ram_depth = 128;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 7;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 127;
defparam ram_block1a18.port_b_logical_ram_depth = 128;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 7;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 127;
defparam ram_block1a17.port_a_logical_ram_depth = 128;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 7;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 127;
defparam ram_block1a17.port_b_logical_ram_depth = 128;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 7;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 127;
defparam ram_block1a31.port_a_logical_ram_depth = 128;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 7;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 127;
defparam ram_block1a31.port_b_logical_ram_depth = 128;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 7;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 127;
defparam ram_block1a30.port_a_logical_ram_depth = 128;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 7;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 127;
defparam ram_block1a30.port_b_logical_ram_depth = 128;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 7;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 127;
defparam ram_block1a29.port_a_logical_ram_depth = 128;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 7;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 127;
defparam ram_block1a29.port_b_logical_ram_depth = 128;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 7;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 127;
defparam ram_block1a28.port_a_logical_ram_depth = 128;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 7;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 127;
defparam ram_block1a28.port_b_logical_ram_depth = 128;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 7;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 127;
defparam ram_block1a27.port_a_logical_ram_depth = 128;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 7;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 127;
defparam ram_block1a27.port_b_logical_ram_depth = 128;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 7;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 127;
defparam ram_block1a26.port_a_logical_ram_depth = 128;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 7;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 127;
defparam ram_block1a26.port_b_logical_ram_depth = 128;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 7;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 127;
defparam ram_block1a25.port_a_logical_ram_depth = 128;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 7;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 127;
defparam ram_block1a25.port_b_logical_ram_depth = 128;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 7;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 127;
defparam ram_block1a24.port_a_logical_ram_depth = 128;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 7;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 127;
defparam ram_block1a24.port_b_logical_ram_depth = 128;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 7;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 127;
defparam ram_block1a23.port_a_logical_ram_depth = 128;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 7;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 127;
defparam ram_block1a23.port_b_logical_ram_depth = 128;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 7;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 127;
defparam ram_block1a22.port_a_logical_ram_depth = 128;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 7;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 127;
defparam ram_block1a22.port_b_logical_ram_depth = 128;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 7;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 127;
defparam ram_block1a20.port_a_logical_ram_depth = 128;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 7;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 127;
defparam ram_block1a20.port_b_logical_ram_depth = 128;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_in_deserializer:Audio_In_Deserializer|altera_up_sync_fifo:Audio_In_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 7;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 127;
defparam ram_block1a19.port_a_logical_ram_depth = 128;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 7;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 127;
defparam ram_block1a19.port_b_logical_ram_depth = 128;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

endmodule

module final_project_soc_cntr_0ab_1 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	clear_read_fifos,
	comb,
	comb1,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_read_fifos;
input 	comb;
input 	comb1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(comb),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFDFD;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_ca7_1 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	altera_reset_synchronizer_int_chain_out,
	clear_read_fifos,
	updown,
	comb,
	comb1,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_read_fifos;
input 	updown;
input 	comb;
input 	comb1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(updown),
	.datad(comb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hDFFD;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_v9b_1 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	altera_reset_synchronizer_int_chain_out,
	clear_read_fifos,
	comb,
	rd_ptr_lsb,
	comb1,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_read_fifos;
input 	comb;
input 	rd_ptr_lsb;
input 	comb1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb1),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_read_fifos),
	.datac(comb),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFDFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_altera_up_audio_out_serializer (
	clk_0,
	done_dac_channel_sync,
	right_channel_fifo_write_space_0,
	right_channel_fifo_write_space_5,
	right_channel_fifo_write_space_2,
	right_channel_fifo_write_space_1,
	left_channel_fifo_write_space_7,
	left_channel_fifo_write_space_6,
	left_channel_fifo_write_space_5,
	left_channel_fifo_write_space_4,
	left_channel_fifo_write_space_3,
	left_channel_fifo_write_space_2,
	left_channel_fifo_write_space_1,
	left_channel_fifo_write_space_0,
	right_channel_fifo_write_space_7,
	right_channel_fifo_write_space_6,
	right_channel_fifo_write_space_4,
	right_channel_fifo_write_space_3,
	serial_audio_out_data1,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	last_test_clk,
	cur_test_clk,
	comb,
	falling_edge,
	src_data_38,
	src_data_39,
	WideOr1,
	mem_used_1,
	nonposted_write_endofpacket,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	done_dac_channel_sync;
output 	right_channel_fifo_write_space_0;
output 	right_channel_fifo_write_space_5;
output 	right_channel_fifo_write_space_2;
output 	right_channel_fifo_write_space_1;
output 	left_channel_fifo_write_space_7;
output 	left_channel_fifo_write_space_6;
output 	left_channel_fifo_write_space_5;
output 	left_channel_fifo_write_space_4;
output 	left_channel_fifo_write_space_3;
output 	left_channel_fifo_write_space_2;
output 	left_channel_fifo_write_space_1;
output 	left_channel_fifo_write_space_0;
output 	right_channel_fifo_write_space_7;
output 	right_channel_fifo_write_space_6;
output 	right_channel_fifo_write_space_4;
output 	right_channel_fifo_write_space_3;
output 	serial_audio_out_data1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	last_test_clk;
input 	cur_test_clk;
input 	comb;
input 	falling_edge;
input 	src_data_38;
input 	src_data_39;
input 	WideOr1;
input 	mem_used_1;
input 	nonposted_write_endofpacket;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \comb~0_combout ;
wire \Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \comb~1_combout ;
wire \Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \comb~2_combout ;
wire \right_channel_fifo_write_space[0]~8_combout ;
wire \right_channel_fifo_write_space[0]~9 ;
wire \right_channel_fifo_write_space[1]~11 ;
wire \right_channel_fifo_write_space[2]~13 ;
wire \right_channel_fifo_write_space[3]~15 ;
wire \right_channel_fifo_write_space[4]~17 ;
wire \right_channel_fifo_write_space[5]~18_combout ;
wire \right_channel_fifo_write_space[2]~12_combout ;
wire \right_channel_fifo_write_space[1]~10_combout ;
wire \left_channel_fifo_write_space[0]~9 ;
wire \left_channel_fifo_write_space[1]~11 ;
wire \left_channel_fifo_write_space[2]~13 ;
wire \left_channel_fifo_write_space[3]~15 ;
wire \left_channel_fifo_write_space[4]~17 ;
wire \left_channel_fifo_write_space[5]~19 ;
wire \left_channel_fifo_write_space[6]~21 ;
wire \left_channel_fifo_write_space[7]~22_combout ;
wire \left_channel_fifo_write_space[6]~20_combout ;
wire \left_channel_fifo_write_space[5]~18_combout ;
wire \left_channel_fifo_write_space[4]~16_combout ;
wire \left_channel_fifo_write_space[3]~14_combout ;
wire \left_channel_fifo_write_space[2]~12_combout ;
wire \left_channel_fifo_write_space[1]~10_combout ;
wire \left_channel_fifo_write_space[0]~8_combout ;
wire \right_channel_fifo_write_space[5]~19 ;
wire \right_channel_fifo_write_space[6]~21 ;
wire \right_channel_fifo_write_space[7]~22_combout ;
wire \right_channel_fifo_write_space[6]~20_combout ;
wire \right_channel_fifo_write_space[4]~16_combout ;
wire \right_channel_fifo_write_space[3]~14_combout ;
wire \always4~0_combout ;
wire \read_left_channel~combout ;
wire \left_channel_was_read~0_combout ;
wire \left_channel_was_read~q ;
wire \read_right_channel~0_combout ;
wire \data_out_shift_reg~36_combout ;
wire \data_out_shift_reg~37_combout ;
wire \data_out_shift_reg~38_combout ;
wire \data_out_shift_reg[0]~q ;
wire \data_out_shift_reg[1]~30_combout ;
wire \data_out_shift_reg[30]~35_combout ;
wire \data_out_shift_reg[30]~39_combout ;
wire \data_out_shift_reg[1]~q ;
wire \data_out_shift_reg[2]~29_combout ;
wire \data_out_shift_reg[2]~q ;
wire \data_out_shift_reg[3]~28_combout ;
wire \data_out_shift_reg[3]~q ;
wire \data_out_shift_reg[4]~27_combout ;
wire \data_out_shift_reg[4]~q ;
wire \data_out_shift_reg[5]~26_combout ;
wire \data_out_shift_reg[5]~q ;
wire \data_out_shift_reg[6]~25_combout ;
wire \data_out_shift_reg[6]~q ;
wire \data_out_shift_reg[7]~24_combout ;
wire \data_out_shift_reg[7]~q ;
wire \data_out_shift_reg[8]~23_combout ;
wire \data_out_shift_reg[8]~q ;
wire \data_out_shift_reg[9]~22_combout ;
wire \data_out_shift_reg[9]~q ;
wire \data_out_shift_reg[10]~21_combout ;
wire \data_out_shift_reg[10]~q ;
wire \data_out_shift_reg[11]~20_combout ;
wire \data_out_shift_reg[11]~q ;
wire \data_out_shift_reg[12]~19_combout ;
wire \data_out_shift_reg[12]~q ;
wire \data_out_shift_reg[13]~18_combout ;
wire \data_out_shift_reg[13]~q ;
wire \data_out_shift_reg[14]~17_combout ;
wire \data_out_shift_reg[14]~q ;
wire \data_out_shift_reg[15]~16_combout ;
wire \data_out_shift_reg[15]~q ;
wire \data_out_shift_reg[16]~15_combout ;
wire \data_out_shift_reg[16]~q ;
wire \data_out_shift_reg[17]~14_combout ;
wire \data_out_shift_reg[17]~q ;
wire \data_out_shift_reg[18]~13_combout ;
wire \data_out_shift_reg[18]~q ;
wire \data_out_shift_reg[19]~12_combout ;
wire \data_out_shift_reg[19]~q ;
wire \data_out_shift_reg[20]~11_combout ;
wire \data_out_shift_reg[20]~q ;
wire \data_out_shift_reg[21]~10_combout ;
wire \data_out_shift_reg[21]~q ;
wire \data_out_shift_reg[22]~9_combout ;
wire \data_out_shift_reg[22]~q ;
wire \data_out_shift_reg[23]~8_combout ;
wire \data_out_shift_reg[23]~q ;
wire \data_out_shift_reg[24]~7_combout ;
wire \data_out_shift_reg[24]~q ;
wire \data_out_shift_reg[25]~6_combout ;
wire \data_out_shift_reg[25]~q ;
wire \data_out_shift_reg[26]~5_combout ;
wire \data_out_shift_reg[26]~q ;
wire \data_out_shift_reg[27]~4_combout ;
wire \data_out_shift_reg[27]~q ;
wire \data_out_shift_reg[28]~3_combout ;
wire \data_out_shift_reg[28]~q ;
wire \data_out_shift_reg[29]~2_combout ;
wire \data_out_shift_reg[29]~q ;
wire \data_out_shift_reg[30]~1_combout ;
wire \data_out_shift_reg[30]~q ;
wire \data_out_shift_reg[31]~0_combout ;
wire \data_out_shift_reg[31]~q ;
wire \serial_audio_out_data~0_combout ;


final_project_soc_altera_up_sync_fifo_3 Audio_Out_Right_Channel_FIFO(
	.clk_0(clk_0),
	.q_b_31(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_30(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_29(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.counter_reg_bit_1(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_6(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.counter_reg_bit_5(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.q_b_28(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_27(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_26(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_25(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_24(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_23(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_22(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_21(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_20(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_19(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_18(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_17(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_16(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_15(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_14(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_13(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_12(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_11(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_10(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_9(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_8(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_7(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_5(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_4(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_3(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_2(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_1(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_0(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_right_channel(\read_right_channel~0_combout ),
	.empty_dff(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(\comb~0_combout ),
	.full_dff(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.comb2(\comb~1_combout ),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.GND_port(GND_port));

final_project_soc_altera_up_sync_fifo_2 Audio_Out_Left_Channel_FIFO(
	.clk_0(clk_0),
	.q_b_31(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_30(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_29(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.counter_reg_bit_1(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_6(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.counter_reg_bit_5(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.q_b_28(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_27(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_26(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_25(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_24(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_23(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_22(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_21(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_20(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_19(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_18(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_17(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_16(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_15(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_14(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_13(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_12(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_11(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_10(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_9(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_8(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_7(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_5(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_4(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_3(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_2(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_1(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_0(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.empty_dff(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.read_left_channel(\read_left_channel~combout ),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(\comb~0_combout ),
	.src_payload(src_payload),
	.full_dff(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.comb2(\comb~2_combout ),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.GND_port(GND_port));

cycloneive_lcell_comb \comb~0 (
	.dataa(src_data_39),
	.datab(WideOr1),
	.datac(nonposted_write_endofpacket),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hFDFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~1 (
	.dataa(src_data_38),
	.datab(\comb~0_combout ),
	.datac(gnd),
	.datad(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'hEEFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~2 (
	.dataa(\comb~0_combout ),
	.datab(gnd),
	.datac(src_data_38),
	.datad(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
defparam \comb~2 .lut_mask = 16'hAFFF;
defparam \comb~2 .sum_lutc_input = "datac";

dffeas \right_channel_fifo_write_space[0] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_0),
	.prn(vcc));
defparam \right_channel_fifo_write_space[0] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[0] .power_up = "low";

dffeas \right_channel_fifo_write_space[5] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_5),
	.prn(vcc));
defparam \right_channel_fifo_write_space[5] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[5] .power_up = "low";

dffeas \right_channel_fifo_write_space[2] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_2),
	.prn(vcc));
defparam \right_channel_fifo_write_space[2] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[2] .power_up = "low";

dffeas \right_channel_fifo_write_space[1] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_1),
	.prn(vcc));
defparam \right_channel_fifo_write_space[1] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[1] .power_up = "low";

dffeas \left_channel_fifo_write_space[7] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_7),
	.prn(vcc));
defparam \left_channel_fifo_write_space[7] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[7] .power_up = "low";

dffeas \left_channel_fifo_write_space[6] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_6),
	.prn(vcc));
defparam \left_channel_fifo_write_space[6] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[6] .power_up = "low";

dffeas \left_channel_fifo_write_space[5] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_5),
	.prn(vcc));
defparam \left_channel_fifo_write_space[5] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[5] .power_up = "low";

dffeas \left_channel_fifo_write_space[4] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_4),
	.prn(vcc));
defparam \left_channel_fifo_write_space[4] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[4] .power_up = "low";

dffeas \left_channel_fifo_write_space[3] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_3),
	.prn(vcc));
defparam \left_channel_fifo_write_space[3] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[3] .power_up = "low";

dffeas \left_channel_fifo_write_space[2] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_2),
	.prn(vcc));
defparam \left_channel_fifo_write_space[2] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[2] .power_up = "low";

dffeas \left_channel_fifo_write_space[1] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_1),
	.prn(vcc));
defparam \left_channel_fifo_write_space[1] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[1] .power_up = "low";

dffeas \left_channel_fifo_write_space[0] (
	.clk(clk_0),
	.d(\left_channel_fifo_write_space[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(left_channel_fifo_write_space_0),
	.prn(vcc));
defparam \left_channel_fifo_write_space[0] .is_wysiwyg = "true";
defparam \left_channel_fifo_write_space[0] .power_up = "low";

dffeas \right_channel_fifo_write_space[7] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_7),
	.prn(vcc));
defparam \right_channel_fifo_write_space[7] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[7] .power_up = "low";

dffeas \right_channel_fifo_write_space[6] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_6),
	.prn(vcc));
defparam \right_channel_fifo_write_space[6] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[6] .power_up = "low";

dffeas \right_channel_fifo_write_space[4] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_4),
	.prn(vcc));
defparam \right_channel_fifo_write_space[4] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[4] .power_up = "low";

dffeas \right_channel_fifo_write_space[3] (
	.clk(clk_0),
	.d(\right_channel_fifo_write_space[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(comb),
	.sload(gnd),
	.ena(vcc),
	.q(right_channel_fifo_write_space_3),
	.prn(vcc));
defparam \right_channel_fifo_write_space[3] .is_wysiwyg = "true";
defparam \right_channel_fifo_write_space[3] .power_up = "low";

dffeas serial_audio_out_data(
	.clk(clk_0),
	.d(\serial_audio_out_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(serial_audio_out_data1),
	.prn(vcc));
defparam serial_audio_out_data.is_wysiwyg = "true";
defparam serial_audio_out_data.power_up = "low";

cycloneive_lcell_comb \right_channel_fifo_write_space[0]~8 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\right_channel_fifo_write_space[0]~8_combout ),
	.cout(\right_channel_fifo_write_space[0]~9 ));
defparam \right_channel_fifo_write_space[0]~8 .lut_mask = 16'hAA55;
defparam \right_channel_fifo_write_space[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \right_channel_fifo_write_space[1]~10 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\right_channel_fifo_write_space[0]~9 ),
	.combout(\right_channel_fifo_write_space[1]~10_combout ),
	.cout(\right_channel_fifo_write_space[1]~11 ));
defparam \right_channel_fifo_write_space[1]~10 .lut_mask = 16'h5AAF;
defparam \right_channel_fifo_write_space[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \right_channel_fifo_write_space[2]~12 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\right_channel_fifo_write_space[1]~11 ),
	.combout(\right_channel_fifo_write_space[2]~12_combout ),
	.cout(\right_channel_fifo_write_space[2]~13 ));
defparam \right_channel_fifo_write_space[2]~12 .lut_mask = 16'h5A5F;
defparam \right_channel_fifo_write_space[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \right_channel_fifo_write_space[3]~14 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\right_channel_fifo_write_space[2]~13 ),
	.combout(\right_channel_fifo_write_space[3]~14_combout ),
	.cout(\right_channel_fifo_write_space[3]~15 ));
defparam \right_channel_fifo_write_space[3]~14 .lut_mask = 16'h5AAF;
defparam \right_channel_fifo_write_space[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \right_channel_fifo_write_space[4]~16 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\right_channel_fifo_write_space[3]~15 ),
	.combout(\right_channel_fifo_write_space[4]~16_combout ),
	.cout(\right_channel_fifo_write_space[4]~17 ));
defparam \right_channel_fifo_write_space[4]~16 .lut_mask = 16'h5A5F;
defparam \right_channel_fifo_write_space[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \right_channel_fifo_write_space[5]~18 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\right_channel_fifo_write_space[4]~17 ),
	.combout(\right_channel_fifo_write_space[5]~18_combout ),
	.cout(\right_channel_fifo_write_space[5]~19 ));
defparam \right_channel_fifo_write_space[5]~18 .lut_mask = 16'h5AAF;
defparam \right_channel_fifo_write_space[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[0]~8 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\left_channel_fifo_write_space[0]~8_combout ),
	.cout(\left_channel_fifo_write_space[0]~9 ));
defparam \left_channel_fifo_write_space[0]~8 .lut_mask = 16'hAA55;
defparam \left_channel_fifo_write_space[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \left_channel_fifo_write_space[1]~10 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\left_channel_fifo_write_space[0]~9 ),
	.combout(\left_channel_fifo_write_space[1]~10_combout ),
	.cout(\left_channel_fifo_write_space[1]~11 ));
defparam \left_channel_fifo_write_space[1]~10 .lut_mask = 16'h5AAF;
defparam \left_channel_fifo_write_space[1]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[2]~12 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\left_channel_fifo_write_space[1]~11 ),
	.combout(\left_channel_fifo_write_space[2]~12_combout ),
	.cout(\left_channel_fifo_write_space[2]~13 ));
defparam \left_channel_fifo_write_space[2]~12 .lut_mask = 16'h5A5F;
defparam \left_channel_fifo_write_space[2]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[3]~14 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\left_channel_fifo_write_space[2]~13 ),
	.combout(\left_channel_fifo_write_space[3]~14_combout ),
	.cout(\left_channel_fifo_write_space[3]~15 ));
defparam \left_channel_fifo_write_space[3]~14 .lut_mask = 16'h5AAF;
defparam \left_channel_fifo_write_space[3]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[4]~16 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\left_channel_fifo_write_space[3]~15 ),
	.combout(\left_channel_fifo_write_space[4]~16_combout ),
	.cout(\left_channel_fifo_write_space[4]~17 ));
defparam \left_channel_fifo_write_space[4]~16 .lut_mask = 16'h5A5F;
defparam \left_channel_fifo_write_space[4]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[5]~18 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\left_channel_fifo_write_space[4]~17 ),
	.combout(\left_channel_fifo_write_space[5]~18_combout ),
	.cout(\left_channel_fifo_write_space[5]~19 ));
defparam \left_channel_fifo_write_space[5]~18 .lut_mask = 16'h5AAF;
defparam \left_channel_fifo_write_space[5]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[6]~20 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\left_channel_fifo_write_space[5]~19 ),
	.combout(\left_channel_fifo_write_space[6]~20_combout ),
	.cout(\left_channel_fifo_write_space[6]~21 ));
defparam \left_channel_fifo_write_space[6]~20 .lut_mask = 16'h5A5F;
defparam \left_channel_fifo_write_space[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \left_channel_fifo_write_space[7]~22 (
	.dataa(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\left_channel_fifo_write_space[6]~21 ),
	.combout(\left_channel_fifo_write_space[7]~22_combout ),
	.cout());
defparam \left_channel_fifo_write_space[7]~22 .lut_mask = 16'h5A5A;
defparam \left_channel_fifo_write_space[7]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \right_channel_fifo_write_space[6]~20 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\right_channel_fifo_write_space[5]~19 ),
	.combout(\right_channel_fifo_write_space[6]~20_combout ),
	.cout(\right_channel_fifo_write_space[6]~21 ));
defparam \right_channel_fifo_write_space[6]~20 .lut_mask = 16'h5A5F;
defparam \right_channel_fifo_write_space[6]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \right_channel_fifo_write_space[7]~22 (
	.dataa(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|full_dff~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\right_channel_fifo_write_space[6]~21 ),
	.combout(\right_channel_fifo_write_space[7]~22_combout ),
	.cout());
defparam \right_channel_fifo_write_space[7]~22 .lut_mask = 16'h5A5A;
defparam \right_channel_fifo_write_space[7]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \always4~0 (
	.dataa(done_dac_channel_sync),
	.datab(gnd),
	.datac(last_test_clk),
	.datad(cur_test_clk),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hAFFA;
defparam \always4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb read_left_channel(
	.dataa(cur_test_clk),
	.datab(\always4~0_combout ),
	.datac(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datad(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.cin(gnd),
	.combout(\read_left_channel~combout ),
	.cout());
defparam read_left_channel.lut_mask = 16'hFFFE;
defparam read_left_channel.sum_lutc_input = "datac";

cycloneive_lcell_comb \left_channel_was_read~0 (
	.dataa(comb),
	.datab(\read_left_channel~combout ),
	.datac(\left_channel_was_read~q ),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\left_channel_was_read~0_combout ),
	.cout());
defparam \left_channel_was_read~0 .lut_mask = 16'hFDFF;
defparam \left_channel_was_read~0 .sum_lutc_input = "datac";

dffeas left_channel_was_read(
	.clk(clk_0),
	.d(\left_channel_was_read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\left_channel_was_read~q ),
	.prn(vcc));
defparam left_channel_was_read.is_wysiwyg = "true";
defparam left_channel_was_read.power_up = "low";

cycloneive_lcell_comb \read_right_channel~0 (
	.dataa(\left_channel_was_read~q ),
	.datab(last_test_clk),
	.datac(done_dac_channel_sync),
	.datad(cur_test_clk),
	.cin(gnd),
	.combout(\read_right_channel~0_combout ),
	.cout());
defparam \read_right_channel~0 .lut_mask = 16'hFEFF;
defparam \read_right_channel~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg~36 (
	.dataa(falling_edge),
	.datab(\data_out_shift_reg[0]~q ),
	.datac(\always4~0_combout ),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~36_combout ),
	.cout());
defparam \data_out_shift_reg~36 .lut_mask = 16'hEFFF;
defparam \data_out_shift_reg~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg~37 (
	.dataa(\data_out_shift_reg~36_combout ),
	.datab(\read_right_channel~0_combout ),
	.datac(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datad(\read_left_channel~combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg~37_combout ),
	.cout());
defparam \data_out_shift_reg~37 .lut_mask = 16'hFEFF;
defparam \data_out_shift_reg~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg~38 (
	.dataa(comb),
	.datab(\data_out_shift_reg~37_combout ),
	.datac(\read_left_channel~combout ),
	.datad(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.cin(gnd),
	.combout(\data_out_shift_reg~38_combout ),
	.cout());
defparam \data_out_shift_reg~38 .lut_mask = 16'hFFFD;
defparam \data_out_shift_reg~38 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[0] (
	.clk(clk_0),
	.d(\data_out_shift_reg~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_out_shift_reg[0]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[0] .is_wysiwyg = "true";
defparam \data_out_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[1]~30 (
	.dataa(\data_out_shift_reg[0]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[1]~30_combout ),
	.cout());
defparam \data_out_shift_reg[1]~30 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[1]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg[30]~35 (
	.dataa(\always4~0_combout ),
	.datab(\read_right_channel~0_combout ),
	.datac(\read_left_channel~combout ),
	.datad(comb),
	.cin(gnd),
	.combout(\data_out_shift_reg[30]~35_combout ),
	.cout());
defparam \data_out_shift_reg[30]~35 .lut_mask = 16'hFFBF;
defparam \data_out_shift_reg[30]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_shift_reg[30]~39 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(falling_edge),
	.datad(\always4~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[30]~39_combout ),
	.cout());
defparam \data_out_shift_reg[30]~39 .lut_mask = 16'hFFDF;
defparam \data_out_shift_reg[30]~39 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[1] (
	.clk(clk_0),
	.d(\data_out_shift_reg[1]~30_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[1]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[1] .is_wysiwyg = "true";
defparam \data_out_shift_reg[1] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[2]~29 (
	.dataa(\data_out_shift_reg[1]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[2]~29_combout ),
	.cout());
defparam \data_out_shift_reg[2]~29 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[2]~29 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[2] (
	.clk(clk_0),
	.d(\data_out_shift_reg[2]~29_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[2]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[2] .is_wysiwyg = "true";
defparam \data_out_shift_reg[2] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[3]~28 (
	.dataa(\data_out_shift_reg[2]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[3]~28_combout ),
	.cout());
defparam \data_out_shift_reg[3]~28 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[3]~28 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[3] (
	.clk(clk_0),
	.d(\data_out_shift_reg[3]~28_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[3]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[3] .is_wysiwyg = "true";
defparam \data_out_shift_reg[3] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[4]~27 (
	.dataa(\data_out_shift_reg[3]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[4]~27_combout ),
	.cout());
defparam \data_out_shift_reg[4]~27 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[4]~27 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[4] (
	.clk(clk_0),
	.d(\data_out_shift_reg[4]~27_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[4]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[4] .is_wysiwyg = "true";
defparam \data_out_shift_reg[4] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[5]~26 (
	.dataa(\data_out_shift_reg[4]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[5]~26_combout ),
	.cout());
defparam \data_out_shift_reg[5]~26 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[5]~26 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[5] (
	.clk(clk_0),
	.d(\data_out_shift_reg[5]~26_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[5]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[5] .is_wysiwyg = "true";
defparam \data_out_shift_reg[5] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[6]~25 (
	.dataa(\data_out_shift_reg[5]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[6]~25_combout ),
	.cout());
defparam \data_out_shift_reg[6]~25 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[6]~25 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[6] (
	.clk(clk_0),
	.d(\data_out_shift_reg[6]~25_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[6]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[6] .is_wysiwyg = "true";
defparam \data_out_shift_reg[6] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[7]~24 (
	.dataa(\data_out_shift_reg[6]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[7]~24_combout ),
	.cout());
defparam \data_out_shift_reg[7]~24 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[7]~24 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[7] (
	.clk(clk_0),
	.d(\data_out_shift_reg[7]~24_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[7]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[7] .is_wysiwyg = "true";
defparam \data_out_shift_reg[7] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[8]~23 (
	.dataa(\data_out_shift_reg[7]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[8]~23_combout ),
	.cout());
defparam \data_out_shift_reg[8]~23 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[8]~23 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[8] (
	.clk(clk_0),
	.d(\data_out_shift_reg[8]~23_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[8]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[8] .is_wysiwyg = "true";
defparam \data_out_shift_reg[8] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[9]~22 (
	.dataa(\data_out_shift_reg[8]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[9]~22_combout ),
	.cout());
defparam \data_out_shift_reg[9]~22 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[9]~22 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[9] (
	.clk(clk_0),
	.d(\data_out_shift_reg[9]~22_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[9]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[9] .is_wysiwyg = "true";
defparam \data_out_shift_reg[9] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[10]~21 (
	.dataa(\data_out_shift_reg[9]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[10]~21_combout ),
	.cout());
defparam \data_out_shift_reg[10]~21 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[10]~21 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[10] (
	.clk(clk_0),
	.d(\data_out_shift_reg[10]~21_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[10]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[10] .is_wysiwyg = "true";
defparam \data_out_shift_reg[10] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[11]~20 (
	.dataa(\data_out_shift_reg[10]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[11]~20_combout ),
	.cout());
defparam \data_out_shift_reg[11]~20 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[11]~20 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[11] (
	.clk(clk_0),
	.d(\data_out_shift_reg[11]~20_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[11]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[11] .is_wysiwyg = "true";
defparam \data_out_shift_reg[11] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[12]~19 (
	.dataa(\data_out_shift_reg[11]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[12]~19_combout ),
	.cout());
defparam \data_out_shift_reg[12]~19 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[12]~19 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[12] (
	.clk(clk_0),
	.d(\data_out_shift_reg[12]~19_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[12]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[12] .is_wysiwyg = "true";
defparam \data_out_shift_reg[12] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[13]~18 (
	.dataa(\data_out_shift_reg[12]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[13]~18_combout ),
	.cout());
defparam \data_out_shift_reg[13]~18 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[13]~18 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[13] (
	.clk(clk_0),
	.d(\data_out_shift_reg[13]~18_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[13]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[13] .is_wysiwyg = "true";
defparam \data_out_shift_reg[13] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[14]~17 (
	.dataa(\data_out_shift_reg[13]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[14]~17_combout ),
	.cout());
defparam \data_out_shift_reg[14]~17 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[14]~17 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[14] (
	.clk(clk_0),
	.d(\data_out_shift_reg[14]~17_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[14]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[14] .is_wysiwyg = "true";
defparam \data_out_shift_reg[14] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[15]~16 (
	.dataa(\data_out_shift_reg[14]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[15]~16_combout ),
	.cout());
defparam \data_out_shift_reg[15]~16 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[15]~16 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[15] (
	.clk(clk_0),
	.d(\data_out_shift_reg[15]~16_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[15]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[15] .is_wysiwyg = "true";
defparam \data_out_shift_reg[15] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[16]~15 (
	.dataa(\data_out_shift_reg[15]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[16]~15_combout ),
	.cout());
defparam \data_out_shift_reg[16]~15 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[16]~15 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[16] (
	.clk(clk_0),
	.d(\data_out_shift_reg[16]~15_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[16]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[16] .is_wysiwyg = "true";
defparam \data_out_shift_reg[16] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[17]~14 (
	.dataa(\data_out_shift_reg[16]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[17]~14_combout ),
	.cout());
defparam \data_out_shift_reg[17]~14 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[17]~14 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[17] (
	.clk(clk_0),
	.d(\data_out_shift_reg[17]~14_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[17]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[17] .is_wysiwyg = "true";
defparam \data_out_shift_reg[17] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[18]~13 (
	.dataa(\data_out_shift_reg[17]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[18]~13_combout ),
	.cout());
defparam \data_out_shift_reg[18]~13 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[18]~13 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[18] (
	.clk(clk_0),
	.d(\data_out_shift_reg[18]~13_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[18]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[18] .is_wysiwyg = "true";
defparam \data_out_shift_reg[18] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[19]~12 (
	.dataa(\data_out_shift_reg[18]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[19]~12_combout ),
	.cout());
defparam \data_out_shift_reg[19]~12 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[19]~12 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[19] (
	.clk(clk_0),
	.d(\data_out_shift_reg[19]~12_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[19]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[19] .is_wysiwyg = "true";
defparam \data_out_shift_reg[19] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[20]~11 (
	.dataa(\data_out_shift_reg[19]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[20]~11_combout ),
	.cout());
defparam \data_out_shift_reg[20]~11 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[20]~11 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[20] (
	.clk(clk_0),
	.d(\data_out_shift_reg[20]~11_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[20]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[20] .is_wysiwyg = "true";
defparam \data_out_shift_reg[20] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[21]~10 (
	.dataa(\data_out_shift_reg[20]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[21]~10_combout ),
	.cout());
defparam \data_out_shift_reg[21]~10 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[21]~10 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[21] (
	.clk(clk_0),
	.d(\data_out_shift_reg[21]~10_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[21]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[21] .is_wysiwyg = "true";
defparam \data_out_shift_reg[21] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[22]~9 (
	.dataa(\data_out_shift_reg[21]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[22]~9_combout ),
	.cout());
defparam \data_out_shift_reg[22]~9 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[22]~9 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[22] (
	.clk(clk_0),
	.d(\data_out_shift_reg[22]~9_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[22]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[22] .is_wysiwyg = "true";
defparam \data_out_shift_reg[22] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[23]~8 (
	.dataa(\data_out_shift_reg[22]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[23]~8_combout ),
	.cout());
defparam \data_out_shift_reg[23]~8 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[23]~8 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[23] (
	.clk(clk_0),
	.d(\data_out_shift_reg[23]~8_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[23]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[23] .is_wysiwyg = "true";
defparam \data_out_shift_reg[23] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[24]~7 (
	.dataa(\data_out_shift_reg[23]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[24]~7_combout ),
	.cout());
defparam \data_out_shift_reg[24]~7 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[24]~7 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[24] (
	.clk(clk_0),
	.d(\data_out_shift_reg[24]~7_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[24]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[24] .is_wysiwyg = "true";
defparam \data_out_shift_reg[24] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[25]~6 (
	.dataa(\data_out_shift_reg[24]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[25]~6_combout ),
	.cout());
defparam \data_out_shift_reg[25]~6 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[25]~6 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[25] (
	.clk(clk_0),
	.d(\data_out_shift_reg[25]~6_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[25]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[25] .is_wysiwyg = "true";
defparam \data_out_shift_reg[25] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[26]~5 (
	.dataa(\data_out_shift_reg[25]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[26]~5_combout ),
	.cout());
defparam \data_out_shift_reg[26]~5 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[26]~5 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[26] (
	.clk(clk_0),
	.d(\data_out_shift_reg[26]~5_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[26]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[26] .is_wysiwyg = "true";
defparam \data_out_shift_reg[26] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[27]~4 (
	.dataa(\data_out_shift_reg[26]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[27]~4_combout ),
	.cout());
defparam \data_out_shift_reg[27]~4 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[27]~4 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[27] (
	.clk(clk_0),
	.d(\data_out_shift_reg[27]~4_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[27]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[27] .is_wysiwyg = "true";
defparam \data_out_shift_reg[27] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[28]~3 (
	.dataa(\data_out_shift_reg[27]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[28]~3_combout ),
	.cout());
defparam \data_out_shift_reg[28]~3 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[28]~3 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[28] (
	.clk(clk_0),
	.d(\data_out_shift_reg[28]~3_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[28]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[28] .is_wysiwyg = "true";
defparam \data_out_shift_reg[28] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[29]~2 (
	.dataa(\data_out_shift_reg[28]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[29]~2_combout ),
	.cout());
defparam \data_out_shift_reg[29]~2 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[29]~2 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[29] (
	.clk(clk_0),
	.d(\data_out_shift_reg[29]~2_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[29]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[29] .is_wysiwyg = "true";
defparam \data_out_shift_reg[29] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[30]~1 (
	.dataa(\data_out_shift_reg[29]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[30]~1_combout ),
	.cout());
defparam \data_out_shift_reg[30]~1 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[30]~1 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[30] (
	.clk(clk_0),
	.d(\data_out_shift_reg[30]~1_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[30]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[30] .is_wysiwyg = "true";
defparam \data_out_shift_reg[30] .power_up = "low";

cycloneive_lcell_comb \data_out_shift_reg[31]~0 (
	.dataa(\data_out_shift_reg[30]~q ),
	.datab(\Audio_Out_Right_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.datac(gnd),
	.datad(\read_right_channel~0_combout ),
	.cin(gnd),
	.combout(\data_out_shift_reg[31]~0_combout ),
	.cout());
defparam \data_out_shift_reg[31]~0 .lut_mask = 16'hAACC;
defparam \data_out_shift_reg[31]~0 .sum_lutc_input = "datac";

dffeas \data_out_shift_reg[31] (
	.clk(clk_0),
	.d(\data_out_shift_reg[31]~0_combout ),
	.asdata(\Audio_Out_Left_Channel_FIFO|Sync_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\data_out_shift_reg[30]~35_combout ),
	.sload(\read_left_channel~combout ),
	.ena(\data_out_shift_reg[30]~39_combout ),
	.q(\data_out_shift_reg[31]~q ),
	.prn(vcc));
defparam \data_out_shift_reg[31] .is_wysiwyg = "true";
defparam \data_out_shift_reg[31] .power_up = "low";

cycloneive_lcell_comb \serial_audio_out_data~0 (
	.dataa(\data_out_shift_reg[31]~q ),
	.datab(altera_reset_synchronizer_int_chain_out),
	.datac(gnd),
	.datad(clear_write_fifos),
	.cin(gnd),
	.combout(\serial_audio_out_data~0_combout ),
	.cout());
defparam \serial_audio_out_data~0 .lut_mask = 16'hEEFF;
defparam \serial_audio_out_data~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_sync_fifo_2 (
	clk_0,
	q_b_31,
	q_b_30,
	q_b_29,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	empty_dff,
	read_left_channel,
	comb,
	src_data_38,
	comb1,
	src_payload,
	full_dff,
	comb2,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
output 	empty_dff;
input 	read_left_channel;
input 	comb;
input 	src_data_38;
input 	comb1;
input 	src_payload;
output 	full_dff;
input 	comb2;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_3 Sync_FIFO(
	.clock(clk_0),
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.empty_dff(empty_dff),
	.read_left_channel(read_left_channel),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.data({src_payload,src_payload1,src_payload2,src_payload3,src_payload4,src_payload5,src_payload6,src_payload7,src_payload8,src_payload9,src_payload10,src_payload11,src_payload12,src_payload13,src_payload14,src_payload15,src_payload16,src_payload17,src_payload18,src_payload19,
src_payload20,src_payload21,src_payload22,src_payload23,src_payload24,src_payload25,src_payload26,src_payload27,src_payload28,src_payload29,src_payload30,src_payload31}),
	.full_dff(full_dff),
	.wrreq(comb2),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_3 (
	clock,
	q,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	empty_dff,
	read_left_channel,
	comb,
	src_data_38,
	comb1,
	data,
	full_dff,
	wrreq,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
output 	empty_dff;
input 	read_left_channel;
input 	comb;
input 	src_data_38;
input 	comb1;
input 	[31:0] data;
output 	full_dff;
input 	wrreq;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_n441_2 auto_generated(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.empty_dff(empty_dff),
	.read_left_channel(read_left_channel),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.full_dff(full_dff),
	.wrreq(wrreq),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_n441_2 (
	clock,
	q,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	empty_dff,
	read_left_channel,
	comb,
	src_data_38,
	comb1,
	data,
	full_dff,
	wrreq,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
output 	empty_dff;
input 	read_left_channel;
input 	comb;
input 	src_data_38;
input 	comb1;
input 	[31:0] data;
output 	full_dff;
input 	wrreq;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_a_dpfifo_as31_2 dpfifo(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.empty_dff1(empty_dff),
	.read_left_channel(read_left_channel),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.full_dff1(full_dff),
	.wreq(wrreq),
	.GND_port(GND_port));

endmodule

module final_project_soc_a_dpfifo_as31_2 (
	clock,
	q,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	empty_dff1,
	read_left_channel,
	comb,
	src_data_38,
	comb1,
	data,
	full_dff1,
	wreq,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
output 	empty_dff1;
input 	read_left_channel;
input 	comb;
input 	src_data_38;
input 	comb1;
input 	[31:0] data;
output 	full_dff1;
input 	wreq;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~2_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \rd_ptr_lsb~3_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_0~2_combout ;
wire \usedw_will_be_0~3_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_2~0_combout ;
wire \_~0_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_will_be_2~2_combout ;
wire \usedw_will_be_2~3_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~1_combout ;
wire \empty_dff~0_combout ;
wire \full_dff~2_combout ;
wire \full_dff~3_combout ;
wire \full_dff~4_combout ;
wire \full_dff~5_combout ;


final_project_soc_cntr_0ab_2 wr_ptr(
	.clock(clock),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.full_dff(full_dff1),
	.GND_port(GND_port));

final_project_soc_cntr_ca7_2 usedw_counter(
	.clock(clock),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_left_channel(read_left_channel),
	.comb(comb),
	.updown(wreq),
	.GND_port(GND_port));

final_project_soc_cntr_v9b_2 rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_left_channel(read_left_channel),
	.comb(comb),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port));

final_project_soc_altsyncram_dh81_2 FIFOram(
	.clock0(clock),
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~3_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(read_left_channel),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(comb),
	.datab(\low_addressa[0]~q ),
	.datac(read_left_channel),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hC5FF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~2 (
	.dataa(clear_write_fifos),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\rd_ptr_lsb~2_combout ),
	.cout());
defparam \rd_ptr_lsb~2 .lut_mask = 16'hFF77;
defparam \rd_ptr_lsb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hDDF5;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hDDF5;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hDDF5;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hDDF5;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datac(\low_addressa[5]~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hDDF5;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datac(\low_addressa[6]~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hDDF5;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(read_left_channel),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~3_combout ),
	.cout());
defparam \rd_ptr_lsb~3 .lut_mask = 16'hFDFD;
defparam \rd_ptr_lsb~3 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

dffeas full_dff(
	.clk(clock),
	.d(\full_dff~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_0~2 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\usedw_will_be_0~2_combout ),
	.cout());
defparam \usedw_will_be_0~2 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(\usedw_will_be_0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_0~3_combout ),
	.cout());
defparam \usedw_will_be_0~3 .lut_mask = 16'hFBFB;
defparam \usedw_will_be_0~3 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(read_left_channel),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(read_left_channel),
	.datab(src_data_38),
	.datac(full_dff1),
	.datad(comb1),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hEFFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~2 (
	.dataa(\usedw_will_be_2~1_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\usedw_will_be_2~2_combout ),
	.cout());
defparam \usedw_will_be_2~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~3 (
	.dataa(comb),
	.datab(\usedw_will_be_2~0_combout ),
	.datac(\_~0_combout ),
	.datad(\usedw_will_be_2~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_2~3_combout ),
	.cout());
defparam \usedw_will_be_2~3 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_2~3 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(comb),
	.datab(\usedw_will_be_1~0_combout ),
	.datac(\usedw_is_2_dff~q ),
	.datad(\_~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(wreq),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(comb),
	.datad(\usedw_will_be_0~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~2 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\full_dff~2_combout ),
	.cout());
defparam \full_dff~2 .lut_mask = 16'hFFFE;
defparam \full_dff~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~3 (
	.dataa(\full_dff~2_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\full_dff~3_combout ),
	.cout());
defparam \full_dff~3 .lut_mask = 16'hFFFE;
defparam \full_dff~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~4 (
	.dataa(full_dff1),
	.datab(wreq),
	.datac(\full_dff~3_combout ),
	.datad(read_left_channel),
	.cin(gnd),
	.combout(\full_dff~4_combout ),
	.cout());
defparam \full_dff~4 .lut_mask = 16'hFBFE;
defparam \full_dff~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(\full_dff~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\full_dff~5_combout ),
	.cout());
defparam \full_dff~5 .lut_mask = 16'hFBFB;
defparam \full_dff~5 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altsyncram_dh81_2 (
	clock0,
	q_b,
	address_a,
	data_a,
	wren_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[6:0] address_a;
input 	[31:0] data_a;
input 	wren_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 7;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 127;
defparam ram_block1a31.port_a_logical_ram_depth = 128;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 7;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 127;
defparam ram_block1a31.port_b_logical_ram_depth = 128;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 7;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 127;
defparam ram_block1a30.port_a_logical_ram_depth = 128;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 7;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 127;
defparam ram_block1a30.port_b_logical_ram_depth = 128;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 7;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 127;
defparam ram_block1a29.port_a_logical_ram_depth = 128;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 7;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 127;
defparam ram_block1a29.port_b_logical_ram_depth = 128;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 7;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 127;
defparam ram_block1a28.port_a_logical_ram_depth = 128;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 7;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 127;
defparam ram_block1a28.port_b_logical_ram_depth = 128;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 7;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 127;
defparam ram_block1a27.port_a_logical_ram_depth = 128;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 7;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 127;
defparam ram_block1a27.port_b_logical_ram_depth = 128;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 7;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 127;
defparam ram_block1a26.port_a_logical_ram_depth = 128;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 7;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 127;
defparam ram_block1a26.port_b_logical_ram_depth = 128;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 7;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 127;
defparam ram_block1a25.port_a_logical_ram_depth = 128;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 7;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 127;
defparam ram_block1a25.port_b_logical_ram_depth = 128;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 7;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 127;
defparam ram_block1a24.port_a_logical_ram_depth = 128;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 7;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 127;
defparam ram_block1a24.port_b_logical_ram_depth = 128;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 7;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 127;
defparam ram_block1a23.port_a_logical_ram_depth = 128;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 7;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 127;
defparam ram_block1a23.port_b_logical_ram_depth = 128;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 7;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 127;
defparam ram_block1a22.port_a_logical_ram_depth = 128;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 7;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 127;
defparam ram_block1a22.port_b_logical_ram_depth = 128;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 7;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 127;
defparam ram_block1a21.port_a_logical_ram_depth = 128;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 7;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 127;
defparam ram_block1a21.port_b_logical_ram_depth = 128;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 7;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 127;
defparam ram_block1a20.port_a_logical_ram_depth = 128;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 7;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 127;
defparam ram_block1a20.port_b_logical_ram_depth = 128;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 7;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 127;
defparam ram_block1a19.port_a_logical_ram_depth = 128;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 7;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 127;
defparam ram_block1a19.port_b_logical_ram_depth = 128;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 7;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 127;
defparam ram_block1a18.port_a_logical_ram_depth = 128;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 7;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 127;
defparam ram_block1a18.port_b_logical_ram_depth = 128;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 7;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 127;
defparam ram_block1a17.port_a_logical_ram_depth = 128;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 7;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 127;
defparam ram_block1a17.port_b_logical_ram_depth = 128;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 7;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 127;
defparam ram_block1a16.port_a_logical_ram_depth = 128;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 7;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 127;
defparam ram_block1a16.port_b_logical_ram_depth = 128;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Left_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module final_project_soc_cntr_0ab_2 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	comb,
	src_data_38,
	comb1,
	full_dff,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	comb;
input 	src_data_38;
input 	comb1;
input 	full_dff;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(comb1),
	.datab(src_data_38),
	.datac(full_dff),
	.datad(comb),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFBF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_ca7_2 (
	clock,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_left_channel,
	comb,
	updown,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_left_channel;
input 	comb;
input 	updown;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(read_left_channel),
	.datad(updown),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hDFFD;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_v9b_2 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_left_channel,
	comb,
	rd_ptr_lsb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_left_channel;
input 	comb;
input 	rd_ptr_lsb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(read_left_channel),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFDFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_altera_up_sync_fifo_3 (
	clk_0,
	q_b_31,
	q_b_30,
	q_b_29,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_right_channel,
	empty_dff,
	comb,
	src_data_38,
	comb1,
	full_dff,
	comb2,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_right_channel;
output 	empty_dff;
input 	comb;
input 	src_data_38;
input 	comb1;
output 	full_dff;
input 	comb2;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_4 Sync_FIFO(
	.clock(clk_0),
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_right_channel(read_right_channel),
	.empty_dff(empty_dff),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.full_dff(full_dff),
	.wrreq(comb2),
	.data({src_payload,src_payload1,src_payload2,src_payload3,src_payload4,src_payload5,src_payload6,src_payload7,src_payload8,src_payload9,src_payload10,src_payload11,src_payload12,src_payload13,src_payload14,src_payload15,src_payload16,src_payload17,src_payload18,src_payload19,
src_payload20,src_payload21,src_payload22,src_payload23,src_payload24,src_payload25,src_payload26,src_payload27,src_payload28,src_payload29,src_payload30,src_payload31}),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_4 (
	clock,
	q,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_right_channel,
	empty_dff,
	comb,
	src_data_38,
	comb1,
	full_dff,
	wrreq,
	data,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_right_channel;
output 	empty_dff;
input 	comb;
input 	src_data_38;
input 	comb1;
output 	full_dff;
input 	wrreq;
input 	[31:0] data;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_n441_3 auto_generated(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_right_channel(read_right_channel),
	.empty_dff(empty_dff),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.full_dff(full_dff),
	.wrreq(wrreq),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.GND_port(GND_port));

endmodule

module final_project_soc_scfifo_n441_3 (
	clock,
	q,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_right_channel,
	empty_dff,
	comb,
	src_data_38,
	comb1,
	full_dff,
	wrreq,
	data,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_right_channel;
output 	empty_dff;
input 	comb;
input 	src_data_38;
input 	comb1;
output 	full_dff;
input 	wrreq;
input 	[31:0] data;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_a_dpfifo_as31_3 dpfifo(
	.clock(clock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_right_channel(read_right_channel),
	.empty_dff1(empty_dff),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.full_dff1(full_dff),
	.wreq(wrreq),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.GND_port(GND_port));

endmodule

module final_project_soc_a_dpfifo_as31_3 (
	clock,
	q,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_right_channel,
	empty_dff1,
	comb,
	src_data_38,
	comb1,
	full_dff1,
	wreq,
	data,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	[31:0] q;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_right_channel;
output 	empty_dff1;
input 	comb;
input 	src_data_38;
input 	comb1;
output 	full_dff1;
input 	wreq;
input 	[31:0] data;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~2_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \low_addressa[5]~5_combout ;
wire \low_addressa[6]~6_combout ;
wire \rd_ptr_lsb~3_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_will_be_0~2_combout ;
wire \usedw_will_be_0~3_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_2~0_combout ;
wire \_~0_combout ;
wire \usedw_will_be_2~1_combout ;
wire \usedw_will_be_2~2_combout ;
wire \usedw_will_be_2~3_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~1_combout ;
wire \empty_dff~0_combout ;
wire \full_dff~2_combout ;
wire \full_dff~3_combout ;
wire \full_dff~4_combout ;
wire \full_dff~5_combout ;


final_project_soc_cntr_0ab_3 wr_ptr(
	.clock(clock),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.comb(comb),
	.src_data_38(src_data_38),
	.comb1(comb1),
	.full_dff(full_dff1),
	.GND_port(GND_port));

final_project_soc_cntr_ca7_3 usedw_counter(
	.clock(clock),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_right_channel(read_right_channel),
	.comb(comb),
	.updown(wreq),
	.GND_port(GND_port));

final_project_soc_cntr_v9b_3 rd_ptr_msb(
	.clock(clock),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clear_write_fifos(clear_write_fifos),
	.read_right_channel(read_right_channel),
	.comb(comb),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port));

final_project_soc_altsyncram_dh81_3 FIFOram(
	.clock0(clock),
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(wreq),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~3_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(read_right_channel),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\low_addressa[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[5]~5 (
	.dataa(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datab(\low_addressa[5]~q ),
	.datac(gnd),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.cout());
defparam \ram_read_address[5]~5 .lut_mask = 16'hAACC;
defparam \ram_read_address[5]~5 .sum_lutc_input = "datac";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\low_addressa[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[6]~6 (
	.dataa(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datab(\low_addressa[6]~q ),
	.datac(gnd),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.cout());
defparam \ram_read_address[6]~6 .lut_mask = 16'hAACC;
defparam \ram_read_address[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(comb),
	.datab(\low_addressa[0]~q ),
	.datac(read_right_channel),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hC5FF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~2 (
	.dataa(clear_write_fifos),
	.datab(\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\rd_ptr_lsb~2_combout ),
	.cout());
defparam \rd_ptr_lsb~2 .lut_mask = 16'hFF77;
defparam \rd_ptr_lsb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hDDF5;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hDDF5;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hDDF5;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hDDF5;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[5]~5 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datac(\low_addressa[5]~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\low_addressa[5]~5_combout ),
	.cout());
defparam \low_addressa[5]~5 .lut_mask = 16'hDDF5;
defparam \low_addressa[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[6]~6 (
	.dataa(comb),
	.datab(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datac(\low_addressa[6]~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\low_addressa[6]~6_combout ),
	.cout());
defparam \low_addressa[6]~6 .lut_mask = 16'hDDF5;
defparam \low_addressa[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(read_right_channel),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~3_combout ),
	.cout());
defparam \rd_ptr_lsb~3 .lut_mask = 16'hFDFD;
defparam \rd_ptr_lsb~3 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

dffeas full_dff(
	.clk(clock),
	.d(\full_dff~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_0~2 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\usedw_will_be_0~2_combout ),
	.cout());
defparam \usedw_will_be_0~2 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_0~3 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(\usedw_will_be_0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_0~3_combout ),
	.cout());
defparam \usedw_will_be_0~3 .lut_mask = 16'hFBFB;
defparam \usedw_will_be_0~3 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\usedw_will_be_0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(wreq),
	.datac(read_right_channel),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~0 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(wreq),
	.datac(\usedw_is_1_dff~q ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\usedw_will_be_2~0_combout ),
	.cout());
defparam \usedw_will_be_2~0 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(read_right_channel),
	.datab(full_dff1),
	.datac(src_data_38),
	.datad(comb1),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hEFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~1 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hEFFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~2 (
	.dataa(\usedw_will_be_2~1_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\usedw_will_be_2~2_combout ),
	.cout());
defparam \usedw_will_be_2~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_2~3 (
	.dataa(comb),
	.datab(\usedw_will_be_2~0_combout ),
	.datac(\_~0_combout ),
	.datad(\usedw_will_be_2~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_2~3_combout ),
	.cout());
defparam \usedw_will_be_2~3 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_2~3 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(comb),
	.datab(\usedw_will_be_1~0_combout ),
	.datac(\usedw_is_2_dff~q ),
	.datad(\_~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFFFD;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(wreq),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(comb),
	.datad(\usedw_will_be_0~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hFF7F;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~2 (
	.dataa(counter_reg_bit_1),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_6),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\full_dff~2_combout ),
	.cout());
defparam \full_dff~2 .lut_mask = 16'hFFFE;
defparam \full_dff~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~3 (
	.dataa(\full_dff~2_combout ),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\full_dff~3_combout ),
	.cout());
defparam \full_dff~3 .lut_mask = 16'hFFFE;
defparam \full_dff~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~4 (
	.dataa(full_dff1),
	.datab(wreq),
	.datac(\full_dff~3_combout ),
	.datad(read_right_channel),
	.cin(gnd),
	.combout(\full_dff~4_combout ),
	.cout());
defparam \full_dff~4 .lut_mask = 16'hFBFE;
defparam \full_dff~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_dff~5 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(\full_dff~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\full_dff~5_combout ),
	.cout());
defparam \full_dff~5 .lut_mask = 16'hFBFB;
defparam \full_dff~5 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altsyncram_dh81_3 (
	clock0,
	q_b,
	address_a,
	wren_a,
	data_a,
	address_b)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[6:0] address_a;
input 	wren_a;
input 	[31:0] data_a;
input 	[6:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 7;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 127;
defparam ram_block1a31.port_a_logical_ram_depth = 128;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 7;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 127;
defparam ram_block1a31.port_b_logical_ram_depth = 128;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 7;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 127;
defparam ram_block1a30.port_a_logical_ram_depth = 128;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 7;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 127;
defparam ram_block1a30.port_b_logical_ram_depth = 128;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 7;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 127;
defparam ram_block1a29.port_a_logical_ram_depth = 128;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 7;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 127;
defparam ram_block1a29.port_b_logical_ram_depth = 128;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 7;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 127;
defparam ram_block1a28.port_a_logical_ram_depth = 128;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 7;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 127;
defparam ram_block1a28.port_b_logical_ram_depth = 128;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 7;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 127;
defparam ram_block1a27.port_a_logical_ram_depth = 128;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 7;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 127;
defparam ram_block1a27.port_b_logical_ram_depth = 128;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 7;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 127;
defparam ram_block1a26.port_a_logical_ram_depth = 128;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 7;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 127;
defparam ram_block1a26.port_b_logical_ram_depth = 128;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 7;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 127;
defparam ram_block1a25.port_a_logical_ram_depth = 128;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 7;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 127;
defparam ram_block1a25.port_b_logical_ram_depth = 128;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 7;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 127;
defparam ram_block1a24.port_a_logical_ram_depth = 128;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 7;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 127;
defparam ram_block1a24.port_b_logical_ram_depth = 128;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 7;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 127;
defparam ram_block1a23.port_a_logical_ram_depth = 128;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 7;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 127;
defparam ram_block1a23.port_b_logical_ram_depth = 128;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 7;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 127;
defparam ram_block1a22.port_a_logical_ram_depth = 128;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 7;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 127;
defparam ram_block1a22.port_b_logical_ram_depth = 128;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 7;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 127;
defparam ram_block1a21.port_a_logical_ram_depth = 128;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 7;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 127;
defparam ram_block1a21.port_b_logical_ram_depth = 128;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 7;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 127;
defparam ram_block1a20.port_a_logical_ram_depth = 128;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 7;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 127;
defparam ram_block1a20.port_b_logical_ram_depth = 128;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 7;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 127;
defparam ram_block1a19.port_a_logical_ram_depth = 128;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 7;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 127;
defparam ram_block1a19.port_b_logical_ram_depth = 128;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 7;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 127;
defparam ram_block1a18.port_a_logical_ram_depth = 128;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 7;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 127;
defparam ram_block1a18.port_b_logical_ram_depth = 128;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 7;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 127;
defparam ram_block1a17.port_a_logical_ram_depth = 128;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 7;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 127;
defparam ram_block1a17.port_b_logical_ram_depth = 128;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 7;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 127;
defparam ram_block1a16.port_a_logical_ram_depth = 128;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 7;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 127;
defparam ram_block1a16.port_b_logical_ram_depth = 128;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 7;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 127;
defparam ram_block1a15.port_a_logical_ram_depth = 128;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 7;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 127;
defparam ram_block1a15.port_b_logical_ram_depth = 128;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 7;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 127;
defparam ram_block1a14.port_a_logical_ram_depth = 128;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 7;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 127;
defparam ram_block1a14.port_b_logical_ram_depth = 128;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 7;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 127;
defparam ram_block1a13.port_a_logical_ram_depth = 128;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 7;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 127;
defparam ram_block1a13.port_b_logical_ram_depth = 128;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 7;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 127;
defparam ram_block1a12.port_a_logical_ram_depth = 128;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 7;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 127;
defparam ram_block1a12.port_b_logical_ram_depth = 128;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 7;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 127;
defparam ram_block1a11.port_a_logical_ram_depth = 128;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 7;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 127;
defparam ram_block1a11.port_b_logical_ram_depth = 128;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 7;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 127;
defparam ram_block1a10.port_a_logical_ram_depth = 128;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 7;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 127;
defparam ram_block1a10.port_b_logical_ram_depth = 128;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_audio:audio|altera_up_audio_out_serializer:Audio_Out_Serializer|altera_up_sync_fifo:Audio_Out_Right_Channel_FIFO|scfifo:Sync_FIFO|scfifo_n441:auto_generated|a_dpfifo_as31:dpfifo|altsyncram_dh81:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module final_project_soc_cntr_0ab_3 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	comb,
	src_data_38,
	comb1,
	full_dff,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	comb;
input 	src_data_38;
input 	comb1;
input 	full_dff;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(src_data_38),
	.datab(comb1),
	.datac(full_dff),
	.datad(comb),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFEF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A5F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_ca7_3 (
	clock,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_6,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_right_channel,
	comb,
	updown,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_6;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_right_channel;
input 	comb;
input 	updown;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~combout ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(read_right_channel),
	.datad(updown),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hDFFD;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout(\counter_comb_bita5~COUT ));
defparam counter_comb_bita5.lut_mask = 16'h5A6F;
defparam counter_comb_bita5.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita6(
	.dataa(counter_reg_bit_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.combout(\counter_comb_bita6~combout ),
	.cout());
defparam counter_comb_bita6.lut_mask = 16'h5A5A;
defparam counter_comb_bita6.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_v9b_3 (
	clock,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	altera_reset_synchronizer_int_chain_out,
	clear_write_fifos,
	read_right_channel,
	comb,
	rd_ptr_lsb,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	altera_reset_synchronizer_int_chain_out;
input 	clear_write_fifos;
input 	read_right_channel;
input 	comb;
input 	rd_ptr_lsb;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~2_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(comb),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(clear_write_fifos),
	.datac(read_right_channel),
	.datad(rd_ptr_lsb),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFDFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_altera_up_clock_edge (
	clk,
	last_test_clk1,
	cur_test_clk1,
	found_edge1,
	test_clk)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	last_test_clk1;
output 	cur_test_clk1;
output 	found_edge1;
input 	test_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas last_test_clk(
	.clk(clk),
	.d(cur_test_clk1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_test_clk1),
	.prn(vcc));
defparam last_test_clk.is_wysiwyg = "true";
defparam last_test_clk.power_up = "low";

dffeas cur_test_clk(
	.clk(clk),
	.d(test_clk),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cur_test_clk1),
	.prn(vcc));
defparam cur_test_clk.is_wysiwyg = "true";
defparam cur_test_clk.power_up = "low";

cycloneive_lcell_comb found_edge(
	.dataa(gnd),
	.datab(gnd),
	.datac(last_test_clk1),
	.datad(cur_test_clk1),
	.cin(gnd),
	.combout(found_edge1),
	.cout());
defparam found_edge.lut_mask = 16'h0FF0;
defparam found_edge.sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_clock_edge_1 (
	clk,
	cur_test_clk1,
	last_test_clk1,
	falling_edge1,
	test_clk)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	cur_test_clk1;
output 	last_test_clk1;
output 	falling_edge1;
input 	test_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas cur_test_clk(
	.clk(clk),
	.d(test_clk),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cur_test_clk1),
	.prn(vcc));
defparam cur_test_clk.is_wysiwyg = "true";
defparam cur_test_clk.power_up = "low";

dffeas last_test_clk(
	.clk(clk),
	.d(cur_test_clk1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_test_clk1),
	.prn(vcc));
defparam last_test_clk.is_wysiwyg = "true";
defparam last_test_clk.power_up = "low";

cycloneive_lcell_comb falling_edge(
	.dataa(cur_test_clk1),
	.datab(gnd),
	.datac(gnd),
	.datad(last_test_clk1),
	.cin(gnd),
	.combout(falling_edge1),
	.cout());
defparam falling_edge.lut_mask = 16'hAAFF;
defparam falling_edge.sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_clock_edge_2 (
	clk,
	last_test_clk1,
	cur_test_clk1,
	test_clk)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	last_test_clk1;
output 	cur_test_clk1;
input 	test_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas last_test_clk(
	.clk(clk),
	.d(cur_test_clk1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_test_clk1),
	.prn(vcc));
defparam last_test_clk.is_wysiwyg = "true";
defparam last_test_clk.power_up = "low";

dffeas cur_test_clk(
	.clk(clk),
	.d(test_clk),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cur_test_clk1),
	.prn(vcc));
defparam cur_test_clk.is_wysiwyg = "true";
defparam cur_test_clk.power_up = "low";

endmodule

module final_project_soc_final_project_soc_audio_config (
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_16,
	readdata_17,
	readdata_8,
	I2C_SCLK,
	saved_grant_1,
	d_write,
	write_accepted,
	src_valid,
	src1_valid,
	saved_grant_0,
	uav_write,
	mem_used_1,
	internal_reset,
	d_writedata_0,
	src_data_32,
	src_data_38,
	src_data_39,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	WideOr1,
	src_data_68,
	waitrequest1,
	Equal2,
	s_serial_transferSTATE_1_PRE_WRITE,
	waitrequest2,
	I2C_SDAT,
	serial_data,
	m0_read,
	readdata_3,
	readdata_4,
	src_payload,
	d_byteenable_2,
	src_payload1,
	readdata_5,
	readdata_7,
	readdata_6,
	d_byteenable_1,
	audio_config_wire_SDAT,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_16;
output 	readdata_17;
output 	readdata_8;
output 	I2C_SCLK;
input 	saved_grant_1;
input 	d_write;
input 	write_accepted;
input 	src_valid;
input 	src1_valid;
input 	saved_grant_0;
input 	uav_write;
input 	mem_used_1;
output 	internal_reset;
input 	d_writedata_0;
input 	src_data_32;
input 	src_data_38;
input 	src_data_39;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	WideOr1;
input 	src_data_68;
output 	waitrequest1;
output 	Equal2;
output 	s_serial_transferSTATE_1_PRE_WRITE;
output 	waitrequest2;
output 	I2C_SDAT;
output 	serial_data;
input 	m0_read;
output 	readdata_3;
output 	readdata_4;
input 	src_payload;
input 	d_byteenable_2;
input 	src_payload1;
output 	readdata_5;
output 	readdata_7;
output 	readdata_6;
input 	d_byteenable_1;
input 	audio_config_wire_SDAT;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \AV_Config_Auto_Init|transfer_data~q ;
wire \AV_Config_Auto_Init|auto_init_complete~q ;
wire \Serial_Bus_Controller|transfer_complete~q ;
wire \AV_Config_Auto_Init|rom_address[4]~q ;
wire \AV_Config_Auto_Init|rom_address[1]~q ;
wire \AV_Config_Auto_Init|rom_address[0]~q ;
wire \AV_Config_Auto_Init|rom_address[2]~q ;
wire \AV_Config_Auto_Init|rom_address[3]~q ;
wire \AV_Config_Auto_Init|rom_address[5]~q ;
wire \Serial_Bus_Controller|shiftreg_data[1]~q ;
wire \Serial_Bus_Controller|shiftreg_data[0]~q ;
wire \Serial_Bus_Controller|shiftreg_data[9]~q ;
wire \Serial_Bus_Controller|shiftreg_data[2]~q ;
wire \Serial_Bus_Controller|shiftreg_data[3]~q ;
wire \Serial_Bus_Controller|shiftreg_data[4]~q ;
wire \Serial_Bus_Controller|shiftreg_data[5]~q ;
wire \AV_Config_Auto_Init|data_out[25]~q ;
wire \Serial_Bus_Controller|shiftreg_data[6]~q ;
wire \AV_Config_Auto_Init|auto_init_error~q ;
wire \Serial_Bus_Controller|shiftreg_data[8]~q ;
wire \Serial_Bus_Controller|shiftreg_data[7]~q ;
wire \AV_Config_Auto_Init|data_out[1]~q ;
wire \external_read_transfer~q ;
wire \AV_Config_Auto_Init|data_out[2]~q ;
wire \AV_Config_Auto_Init|data_out[3]~q ;
wire \AV_Config_Auto_Init|data_out[4]~q ;
wire \AV_Config_Auto_Init|data_out[5]~q ;
wire \AV_Config_Auto_Init|data_out[6]~q ;
wire \AV_Config_Auto_Init|data_out[10]~q ;
wire \data_reg[8]~q ;
wire \AV_Config_Auto_Init|data_out[8]~q ;
wire \AV_Config_Auto_Init|data_out[7]~q ;
wire \AV_Config_Auto_Init|data_out[17]~q ;
wire \AV_Config_Auto_Init|data_out[16]~q ;
wire \AV_Config_Auto_Init|data_out[15]~q ;
wire \AV_Config_Auto_Init|data_out[14]~q ;
wire \AV_Config_Auto_Init|data_out[13]~q ;
wire \AV_Config_Auto_Init|data_out[12]~q ;
wire \AV_Config_Auto_Init|data_out[11]~q ;
wire \Serial_Bus_Controller|shiftreg_mask~2_combout ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~0_combout ;
wire \Serial_Bus_Controller|shiftreg_data[18]~q ;
wire \device_for_transfer[1]~q ;
wire \device_for_transfer[0]~q ;
wire \Serial_Bus_Controller|shiftreg_data[10]~q ;
wire \data_reg[0]~q ;
wire \Equal5~0_combout ;
wire \data_reg[1]~q ;
wire \data_reg[2]~q ;
wire \data_reg[3]~q ;
wire \data_reg[4]~q ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~3_combout ;
wire \device_for_transfer~0_combout ;
wire \device_for_transfer[0]~1_combout ;
wire \device_for_transfer~2_combout ;
wire \AV_Config_Auto_Init|data_out[24]~q ;
wire \data_reg[5]~q ;
wire \address_for_transfer[0]~q ;
wire \data_reg[7]~q ;
wire \data_reg[6]~q ;
wire \data_reg[0]~2_combout ;
wire \address_for_transfer[7]~q ;
wire \address_for_transfer[6]~q ;
wire \external_read_transfer~0_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[2]~45_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[3]~52_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[4]~combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[5]~57_combout ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Audio_ROM|WideOr0~0_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[6]~58_combout ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~15_combout ;
wire \address_for_transfer~0_combout ;
wire \always3~0_combout ;
wire \data_reg~3_combout ;
wire \data_reg~4_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[8]~61_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[7]~67_combout ;
wire \address_for_transfer~1_combout ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~20_combout ;
wire \address_for_transfer[5]~q ;
wire \address_for_transfer~2_combout ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~22_combout ;
wire \address_for_transfer[4]~q ;
wire \address_for_transfer~3_combout ;
wire \Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~25_combout ;
wire \address_for_transfer[3]~q ;
wire \address_for_transfer~4_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[14]~72_combout ;
wire \address_for_transfer[2]~q ;
wire \address_for_transfer~5_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[13]~77_combout ;
wire \address_for_transfer[1]~q ;
wire \address_for_transfer~6_combout ;
wire \address_for_transfer~7_combout ;
wire \data_reg[0]~5_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[11]~32_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[1]~34_combout ;
wire \Auto_Init_OB_Devices_ROM|rom_data[12]~36_combout ;
wire \ack~0_combout ;
wire \readdata~0_combout ;
wire \address_reg~0_combout ;
wire \address_reg[4]~1_combout ;
wire \address_reg[4]~2_combout ;
wire \address_reg[0]~q ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \control_reg~3_combout ;
wire \address_reg[1]~q ;
wire \internal_reset~3_combout ;
wire \s_serial_transfer~12_combout ;
wire \Selector2~0_combout ;
wire \s_serial_transfer.STATE_5_READ_TRANSFER~q ;
wire \Selector3~0_combout ;
wire \control_reg[17]~0_combout ;
wire \control_reg[17]~1_combout ;
wire \control_reg[17]~2_combout ;
wire \control_reg[16]~q ;
wire \control_reg[17]~q ;
wire \Selector3~1_combout ;
wire \s_serial_transfer.STATE_6_POST_READ~q ;
wire \ns_serial_transfer~2_combout ;
wire \s_serial_transfer~18_combout ;
wire \s_serial_transfer~19_combout ;
wire \Selector1~0_combout ;
wire \s_serial_transfer.STATE_2_WRITE_TRANSFER~q ;
wire \s_serial_transfer~21_combout ;
wire \s_serial_transfer.STATE_3_POST_WRITE~q ;
wire \s_serial_transfer~20_combout ;
wire \s_serial_transfer.STATE_0_IDLE~q ;
wire \s_serial_transfer~13_combout ;
wire \s_serial_transfer~14_combout ;
wire \s_serial_transfer~17_combout ;
wire \s_serial_transfer.STATE_4_PRE_READ~q ;
wire \start_external_transfer~0_combout ;
wire \start_external_transfer~q ;
wire \readdata~3_combout ;
wire \control_reg[2]~4_combout ;
wire \control_reg[2]~5_combout ;
wire \control_reg[1]~q ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \control_reg~6_combout ;
wire \address_reg[2]~q ;
wire \control_reg[2]~q ;
wire \readdata~8_combout ;
wire \readdata~9_combout ;
wire \readdata~14_combout ;
wire \readdata[3]~12_combout ;
wire \readdata~16_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;
wire \internal_reset~4_combout ;
wire \waitrequest~0_combout ;
wire \s_serial_transfer~15_combout ;
wire \s_serial_transfer~16_combout ;
wire \readdata[3]~10_combout ;
wire \address_reg~3_combout ;
wire \address_reg[3]~q ;
wire \readdata~11_combout ;
wire \address_reg~4_combout ;
wire \address_reg[4]~q ;
wire \readdata~13_combout ;
wire \address_reg~5_combout ;
wire \address_reg[5]~q ;
wire \readdata~15_combout ;
wire \address_reg~6_combout ;
wire \address_reg[7]~q ;
wire \readdata~20_combout ;
wire \address_reg~7_combout ;
wire \address_reg[6]~q ;
wire \readdata~21_combout ;


final_project_soc_altera_up_av_config_serial_bus_controller Serial_Bus_Controller(
	.transfer_data(\AV_Config_Auto_Init|transfer_data~q ),
	.auto_init_complete(\AV_Config_Auto_Init|auto_init_complete~q ),
	.transfer_complete1(\Serial_Bus_Controller|transfer_complete~q ),
	.shiftreg_data_1(\Serial_Bus_Controller|shiftreg_data[1]~q ),
	.shiftreg_data_0(\Serial_Bus_Controller|shiftreg_data[0]~q ),
	.shiftreg_data_9(\Serial_Bus_Controller|shiftreg_data[9]~q ),
	.shiftreg_data_2(\Serial_Bus_Controller|shiftreg_data[2]~q ),
	.shiftreg_data_3(\Serial_Bus_Controller|shiftreg_data[3]~q ),
	.shiftreg_data_4(\Serial_Bus_Controller|shiftreg_data[4]~q ),
	.shiftreg_data_5(\Serial_Bus_Controller|shiftreg_data[5]~q ),
	.data_out_25(\AV_Config_Auto_Init|data_out[25]~q ),
	.shiftreg_data_6(\Serial_Bus_Controller|shiftreg_data[6]~q ),
	.shiftreg_data_8(\Serial_Bus_Controller|shiftreg_data[8]~q ),
	.shiftreg_data_7(\Serial_Bus_Controller|shiftreg_data[7]~q ),
	.data_out_1(\AV_Config_Auto_Init|data_out[1]~q ),
	.external_read_transfer(\external_read_transfer~q ),
	.data_out_2(\AV_Config_Auto_Init|data_out[2]~q ),
	.data_out_3(\AV_Config_Auto_Init|data_out[3]~q ),
	.data_out_4(\AV_Config_Auto_Init|data_out[4]~q ),
	.data_out_5(\AV_Config_Auto_Init|data_out[5]~q ),
	.data_out_6(\AV_Config_Auto_Init|data_out[6]~q ),
	.data_out_10(\AV_Config_Auto_Init|data_out[10]~q ),
	.data_reg_8(\data_reg[8]~q ),
	.data_out_8(\AV_Config_Auto_Init|data_out[8]~q ),
	.data_out_7(\AV_Config_Auto_Init|data_out[7]~q ),
	.data_out_17(\AV_Config_Auto_Init|data_out[17]~q ),
	.data_out_16(\AV_Config_Auto_Init|data_out[16]~q ),
	.data_out_15(\AV_Config_Auto_Init|data_out[15]~q ),
	.data_out_14(\AV_Config_Auto_Init|data_out[14]~q ),
	.data_out_13(\AV_Config_Auto_Init|data_out[13]~q ),
	.data_out_12(\AV_Config_Auto_Init|data_out[12]~q ),
	.data_out_11(\AV_Config_Auto_Init|data_out[11]~q ),
	.serial_clk(I2C_SCLK),
	.internal_reset(internal_reset),
	.internal_reset1(\internal_reset~3_combout ),
	.r_sync_rst(r_sync_rst),
	.start_external_transfer(\start_external_transfer~q ),
	.shiftreg_mask(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.serial_data(I2C_SDAT),
	.serial_data1(serial_data),
	.shiftreg_data_18(\Serial_Bus_Controller|shiftreg_data[18]~q ),
	.ack(\ack~0_combout ),
	.device_for_transfer_1(\device_for_transfer[1]~q ),
	.device_for_transfer_0(\device_for_transfer[0]~q ),
	.shiftreg_data_10(\Serial_Bus_Controller|shiftreg_data[10]~q ),
	.data_reg_0(\data_reg[0]~q ),
	.Equal5(\Equal5~0_combout ),
	.data_reg_1(\data_reg[1]~q ),
	.data_reg_2(\data_reg[2]~q ),
	.data_reg_3(\data_reg[3]~q ),
	.data_reg_4(\data_reg[4]~q ),
	.data_out_24(\AV_Config_Auto_Init|data_out[24]~q ),
	.data_reg_5(\data_reg[5]~q ),
	.address_for_transfer_0(\address_for_transfer[0]~q ),
	.data_reg_7(\data_reg[7]~q ),
	.data_reg_6(\data_reg[6]~q ),
	.address_for_transfer_7(\address_for_transfer[7]~q ),
	.address_for_transfer_6(\address_for_transfer[6]~q ),
	.address_for_transfer_5(\address_for_transfer[5]~q ),
	.address_for_transfer_4(\address_for_transfer[4]~q ),
	.address_for_transfer_3(\address_for_transfer[3]~q ),
	.address_for_transfer_2(\address_for_transfer[2]~q ),
	.address_for_transfer_1(\address_for_transfer[1]~q ),
	.audio_config_wire_SDAT(audio_config_wire_SDAT),
	.clk_clk(clk_clk));

final_project_soc_altera_up_av_config_auto_init_ob_de2_115 Auto_Init_OB_Devices_ROM(
	.rom_address_4(\AV_Config_Auto_Init|rom_address[4]~q ),
	.rom_address_1(\AV_Config_Auto_Init|rom_address[1]~q ),
	.rom_address_0(\AV_Config_Auto_Init|rom_address[0]~q ),
	.rom_address_2(\AV_Config_Auto_Init|rom_address[2]~q ),
	.rom_address_3(\AV_Config_Auto_Init|rom_address[3]~q ),
	.rom_address_5(\AV_Config_Auto_Init|rom_address[5]~q ),
	.Ram0(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~0_combout ),
	.Ram01(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~3_combout ),
	.rom_data_2(\Auto_Init_OB_Devices_ROM|rom_data[2]~45_combout ),
	.rom_data_3(\Auto_Init_OB_Devices_ROM|rom_data[3]~52_combout ),
	.rom_data_4(\Auto_Init_OB_Devices_ROM|rom_data[4]~combout ),
	.rom_data_5(\Auto_Init_OB_Devices_ROM|rom_data[5]~57_combout ),
	.WideOr0(\Auto_Init_OB_Devices_ROM|Auto_Init_Audio_ROM|WideOr0~0_combout ),
	.rom_data_6(\Auto_Init_OB_Devices_ROM|rom_data[6]~58_combout ),
	.Ram02(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~15_combout ),
	.rom_data_8(\Auto_Init_OB_Devices_ROM|rom_data[8]~61_combout ),
	.rom_data_7(\Auto_Init_OB_Devices_ROM|rom_data[7]~67_combout ),
	.Ram03(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~20_combout ),
	.Ram04(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~22_combout ),
	.Ram05(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~25_combout ),
	.rom_data_14(\Auto_Init_OB_Devices_ROM|rom_data[14]~72_combout ),
	.rom_data_13(\Auto_Init_OB_Devices_ROM|rom_data[13]~77_combout ),
	.rom_data_11(\Auto_Init_OB_Devices_ROM|rom_data[11]~32_combout ),
	.rom_data_1(\Auto_Init_OB_Devices_ROM|rom_data[1]~34_combout ),
	.rom_data_12(\Auto_Init_OB_Devices_ROM|rom_data[12]~36_combout ));

final_project_soc_altera_up_av_config_auto_init AV_Config_Auto_Init(
	.transfer_data1(\AV_Config_Auto_Init|transfer_data~q ),
	.auto_init_complete1(\AV_Config_Auto_Init|auto_init_complete~q ),
	.transfer_complete(\Serial_Bus_Controller|transfer_complete~q ),
	.rom_address_4(\AV_Config_Auto_Init|rom_address[4]~q ),
	.rom_address_1(\AV_Config_Auto_Init|rom_address[1]~q ),
	.rom_address_0(\AV_Config_Auto_Init|rom_address[0]~q ),
	.rom_address_2(\AV_Config_Auto_Init|rom_address[2]~q ),
	.rom_address_3(\AV_Config_Auto_Init|rom_address[3]~q ),
	.rom_address_5(\AV_Config_Auto_Init|rom_address[5]~q ),
	.data_out_25(\AV_Config_Auto_Init|data_out[25]~q ),
	.auto_init_error1(\AV_Config_Auto_Init|auto_init_error~q ),
	.data_out_1(\AV_Config_Auto_Init|data_out[1]~q ),
	.data_out_2(\AV_Config_Auto_Init|data_out[2]~q ),
	.data_out_3(\AV_Config_Auto_Init|data_out[3]~q ),
	.data_out_4(\AV_Config_Auto_Init|data_out[4]~q ),
	.data_out_5(\AV_Config_Auto_Init|data_out[5]~q ),
	.data_out_6(\AV_Config_Auto_Init|data_out[6]~q ),
	.data_out_10(\AV_Config_Auto_Init|data_out[10]~q ),
	.data_out_8(\AV_Config_Auto_Init|data_out[8]~q ),
	.data_out_7(\AV_Config_Auto_Init|data_out[7]~q ),
	.data_out_17(\AV_Config_Auto_Init|data_out[17]~q ),
	.data_out_16(\AV_Config_Auto_Init|data_out[16]~q ),
	.data_out_15(\AV_Config_Auto_Init|data_out[15]~q ),
	.data_out_14(\AV_Config_Auto_Init|data_out[14]~q ),
	.data_out_13(\AV_Config_Auto_Init|data_out[13]~q ),
	.data_out_12(\AV_Config_Auto_Init|data_out[12]~q ),
	.data_out_11(\AV_Config_Auto_Init|data_out[11]~q ),
	.shiftreg_mask(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.Ram0(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~0_combout ),
	.ack(\ack~0_combout ),
	.Ram01(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~3_combout ),
	.data_out_24(\AV_Config_Auto_Init|data_out[24]~q ),
	.rom_data_2(\Auto_Init_OB_Devices_ROM|rom_data[2]~45_combout ),
	.rom_data_3(\Auto_Init_OB_Devices_ROM|rom_data[3]~52_combout ),
	.rom_data_4(\Auto_Init_OB_Devices_ROM|rom_data[4]~combout ),
	.rom_data_5(\Auto_Init_OB_Devices_ROM|rom_data[5]~57_combout ),
	.WideOr0(\Auto_Init_OB_Devices_ROM|Auto_Init_Audio_ROM|WideOr0~0_combout ),
	.rom_data_6(\Auto_Init_OB_Devices_ROM|rom_data[6]~58_combout ),
	.Ram02(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~15_combout ),
	.rom_data_8(\Auto_Init_OB_Devices_ROM|rom_data[8]~61_combout ),
	.rom_data_7(\Auto_Init_OB_Devices_ROM|rom_data[7]~67_combout ),
	.Ram03(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~20_combout ),
	.Ram04(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~22_combout ),
	.Ram05(\Auto_Init_OB_Devices_ROM|Auto_Init_Video_ROM|Ram0~25_combout ),
	.rom_data_14(\Auto_Init_OB_Devices_ROM|rom_data[14]~72_combout ),
	.rom_data_13(\Auto_Init_OB_Devices_ROM|rom_data[13]~77_combout ),
	.rom_data_11(\Auto_Init_OB_Devices_ROM|rom_data[11]~32_combout ),
	.rom_data_1(\Auto_Init_OB_Devices_ROM|rom_data[1]~34_combout ),
	.rom_data_12(\Auto_Init_OB_Devices_ROM|rom_data[12]~36_combout ),
	.clk_clk(clk_clk));

dffeas external_read_transfer(
	.clk(clk_clk),
	.d(\external_read_transfer~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\external_read_transfer~q ),
	.prn(vcc));
defparam external_read_transfer.is_wysiwyg = "true";
defparam external_read_transfer.power_up = "low";

dffeas \data_reg[8] (
	.clk(clk_clk),
	.d(\data_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[8]~q ),
	.prn(vcc));
defparam \data_reg[8] .is_wysiwyg = "true";
defparam \data_reg[8] .power_up = "low";

dffeas \device_for_transfer[1] (
	.clk(clk_clk),
	.d(\device_for_transfer~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\device_for_transfer[0]~1_combout ),
	.q(\device_for_transfer[1]~q ),
	.prn(vcc));
defparam \device_for_transfer[1] .is_wysiwyg = "true";
defparam \device_for_transfer[1] .power_up = "low";

dffeas \device_for_transfer[0] (
	.clk(clk_clk),
	.d(\device_for_transfer~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\device_for_transfer[0]~1_combout ),
	.q(\device_for_transfer[0]~q ),
	.prn(vcc));
defparam \device_for_transfer[0] .is_wysiwyg = "true";
defparam \device_for_transfer[0] .power_up = "low";

dffeas \data_reg[0] (
	.clk(clk_clk),
	.d(\address_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[0]~q ),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

cycloneive_lcell_comb \Equal5~0 (
	.dataa(\device_for_transfer[1]~q ),
	.datab(\device_for_transfer[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'hEEEE;
defparam \Equal5~0 .sum_lutc_input = "datac";

dffeas \data_reg[1] (
	.clk(clk_clk),
	.d(\control_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[1]~q ),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

dffeas \data_reg[2] (
	.clk(clk_clk),
	.d(\control_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[2]~q ),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

dffeas \data_reg[3] (
	.clk(clk_clk),
	.d(\address_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[3]~q ),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

dffeas \data_reg[4] (
	.clk(clk_clk),
	.d(\address_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[4]~q ),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

cycloneive_lcell_comb \device_for_transfer~0 (
	.dataa(\control_reg[17]~q ),
	.datab(internal_reset),
	.datac(\internal_reset~3_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\device_for_transfer~0_combout ),
	.cout());
defparam \device_for_transfer~0 .lut_mask = 16'hBFFF;
defparam \device_for_transfer~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \device_for_transfer[0]~1 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(\Serial_Bus_Controller|transfer_complete~q ),
	.datac(s_serial_transferSTATE_1_PRE_WRITE),
	.datad(\s_serial_transfer.STATE_4_PRE_READ~q ),
	.cin(gnd),
	.combout(\device_for_transfer[0]~1_combout ),
	.cout());
defparam \device_for_transfer[0]~1 .lut_mask = 16'hFFFB;
defparam \device_for_transfer[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \device_for_transfer~2 (
	.dataa(\control_reg[16]~q ),
	.datab(internal_reset),
	.datac(\internal_reset~3_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\device_for_transfer~2_combout ),
	.cout());
defparam \device_for_transfer~2 .lut_mask = 16'hBFFF;
defparam \device_for_transfer~2 .sum_lutc_input = "datac";

dffeas \data_reg[5] (
	.clk(clk_clk),
	.d(\address_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[5]~q ),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

dffeas \address_for_transfer[0] (
	.clk(clk_clk),
	.d(\address_for_transfer~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[0]~q ),
	.prn(vcc));
defparam \address_for_transfer[0] .is_wysiwyg = "true";
defparam \address_for_transfer[0] .power_up = "low";

dffeas \data_reg[7] (
	.clk(clk_clk),
	.d(\address_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[7]~q ),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

dffeas \data_reg[6] (
	.clk(clk_clk),
	.d(\address_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_reg[0]~2_combout ),
	.q(\data_reg[6]~q ),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

cycloneive_lcell_comb \data_reg[0]~2 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(internal_reset),
	.datac(waitrequest1),
	.datad(\data_reg[0]~5_combout ),
	.cin(gnd),
	.combout(\data_reg[0]~2_combout ),
	.cout());
defparam \data_reg[0]~2 .lut_mask = 16'hEFFF;
defparam \data_reg[0]~2 .sum_lutc_input = "datac";

dffeas \address_for_transfer[7] (
	.clk(clk_clk),
	.d(\address_for_transfer~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[7]~q ),
	.prn(vcc));
defparam \address_for_transfer[7] .is_wysiwyg = "true";
defparam \address_for_transfer[7] .power_up = "low";

dffeas \address_for_transfer[6] (
	.clk(clk_clk),
	.d(\address_for_transfer~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[6]~q ),
	.prn(vcc));
defparam \address_for_transfer[6] .is_wysiwyg = "true";
defparam \address_for_transfer[6] .power_up = "low";

cycloneive_lcell_comb \external_read_transfer~0 (
	.dataa(\Serial_Bus_Controller|transfer_complete~q ),
	.datab(s_serial_transferSTATE_1_PRE_WRITE),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\external_read_transfer~0_combout ),
	.cout());
defparam \external_read_transfer~0 .lut_mask = 16'h7777;
defparam \external_read_transfer~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_for_transfer~0 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~0_combout ),
	.cout());
defparam \address_for_transfer~0 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always3~0 (
	.dataa(internal_reset),
	.datab(s_serial_transferSTATE_1_PRE_WRITE),
	.datac(Equal2),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hEFFF;
defparam \always3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~3 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(saved_grant_1),
	.datad(d_byteenable_1),
	.cin(gnd),
	.combout(\data_reg~3_combout ),
	.cout());
defparam \data_reg~3 .lut_mask = 16'hFFFE;
defparam \data_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg~4 (
	.dataa(d_writedata_8),
	.datab(\data_reg[8]~q ),
	.datac(\always3~0_combout ),
	.datad(\data_reg~3_combout ),
	.cin(gnd),
	.combout(\data_reg~4_combout ),
	.cout());
defparam \data_reg~4 .lut_mask = 16'hEFFE;
defparam \data_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_for_transfer~1 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~1_combout ),
	.cout());
defparam \address_for_transfer~1 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~1 .sum_lutc_input = "datac";

dffeas \address_for_transfer[5] (
	.clk(clk_clk),
	.d(\address_for_transfer~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[5]~q ),
	.prn(vcc));
defparam \address_for_transfer[5] .is_wysiwyg = "true";
defparam \address_for_transfer[5] .power_up = "low";

cycloneive_lcell_comb \address_for_transfer~2 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~2_combout ),
	.cout());
defparam \address_for_transfer~2 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~2 .sum_lutc_input = "datac";

dffeas \address_for_transfer[4] (
	.clk(clk_clk),
	.d(\address_for_transfer~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[4]~q ),
	.prn(vcc));
defparam \address_for_transfer[4] .is_wysiwyg = "true";
defparam \address_for_transfer[4] .power_up = "low";

cycloneive_lcell_comb \address_for_transfer~3 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~3_combout ),
	.cout());
defparam \address_for_transfer~3 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~3 .sum_lutc_input = "datac";

dffeas \address_for_transfer[3] (
	.clk(clk_clk),
	.d(\address_for_transfer~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[3]~q ),
	.prn(vcc));
defparam \address_for_transfer[3] .is_wysiwyg = "true";
defparam \address_for_transfer[3] .power_up = "low";

cycloneive_lcell_comb \address_for_transfer~4 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~4_combout ),
	.cout());
defparam \address_for_transfer~4 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~4 .sum_lutc_input = "datac";

dffeas \address_for_transfer[2] (
	.clk(clk_clk),
	.d(\address_for_transfer~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[2]~q ),
	.prn(vcc));
defparam \address_for_transfer[2] .is_wysiwyg = "true";
defparam \address_for_transfer[2] .power_up = "low";

cycloneive_lcell_comb \address_for_transfer~5 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~5_combout ),
	.cout());
defparam \address_for_transfer~5 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~5 .sum_lutc_input = "datac";

dffeas \address_for_transfer[1] (
	.clk(clk_clk),
	.d(\address_for_transfer~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\address_for_transfer[1]~q ),
	.prn(vcc));
defparam \address_for_transfer[1] .is_wysiwyg = "true";
defparam \address_for_transfer[1] .power_up = "low";

cycloneive_lcell_comb \address_for_transfer~6 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~6_combout ),
	.cout());
defparam \address_for_transfer~6 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_for_transfer~7 (
	.dataa(\s_serial_transfer~12_combout ),
	.datab(\address_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_for_transfer~7_combout ),
	.cout());
defparam \address_for_transfer~7 .lut_mask = 16'hEEEE;
defparam \address_for_transfer~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_reg[0]~5 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(src_data_32),
	.datad(s_serial_transferSTATE_1_PRE_WRITE),
	.cin(gnd),
	.combout(\data_reg[0]~5_combout ),
	.cout());
defparam \data_reg[0]~5 .lut_mask = 16'h7FFF;
defparam \data_reg[0]~5 .sum_lutc_input = "datac";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

cycloneive_lcell_comb \internal_reset~2 (
	.dataa(saved_grant_1),
	.datab(src_valid),
	.datac(src1_valid),
	.datad(\internal_reset~4_combout ),
	.cin(gnd),
	.combout(internal_reset),
	.cout());
defparam \internal_reset~2 .lut_mask = 16'hFFFE;
defparam \internal_reset~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \waitrequest~1 (
	.dataa(WideOr1),
	.datab(src_data_68),
	.datac(\waitrequest~0_combout ),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(waitrequest1),
	.cout());
defparam \waitrequest~1 .lut_mask = 16'hFEFF;
defparam \waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEEEE;
defparam \Equal2~0 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_1_PRE_WRITE (
	.clk(clk_clk),
	.d(\s_serial_transfer~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(s_serial_transferSTATE_1_PRE_WRITE),
	.prn(vcc));
defparam \s_serial_transfer.STATE_1_PRE_WRITE .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_1_PRE_WRITE .power_up = "low";

cycloneive_lcell_comb waitrequest(
	.dataa(waitrequest1),
	.datab(internal_reset),
	.datac(Equal2),
	.datad(s_serial_transferSTATE_1_PRE_WRITE),
	.cin(gnd),
	.combout(waitrequest2),
	.cout());
defparam waitrequest.lut_mask = 16'hFEFF;
defparam waitrequest.sum_lutc_input = "datac";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata[3]~12_combout ),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

cycloneive_lcell_comb \ack~0 (
	.dataa(\Serial_Bus_Controller|shiftreg_data[18]~q ),
	.datab(\Serial_Bus_Controller|shiftreg_data[0]~q ),
	.datac(\Serial_Bus_Controller|shiftreg_data[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ack~0_combout ),
	.cout());
defparam \ack~0 .lut_mask = 16'hFEFE;
defparam \ack~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~0 (
	.dataa(src_data_38),
	.datab(\Serial_Bus_Controller|shiftreg_data[1]~q ),
	.datac(\ack~0_combout ),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hFAFC;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~0 (
	.dataa(saved_grant_0),
	.datab(d_writedata_0),
	.datac(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg~0_combout ),
	.cout());
defparam \address_reg~0 .lut_mask = 16'hEFEF;
defparam \address_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg[4]~1 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(src_data_32),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg[4]~1_combout ),
	.cout());
defparam \address_reg[4]~1 .lut_mask = 16'hBFBF;
defparam \address_reg[4]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg[4]~2 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(internal_reset),
	.datac(waitrequest2),
	.datad(\address_reg[4]~1_combout ),
	.cin(gnd),
	.combout(\address_reg[4]~2_combout ),
	.cout());
defparam \address_reg[4]~2 .lut_mask = 16'hEFFF;
defparam \address_reg[4]~2 .sum_lutc_input = "datac";

dffeas \address_reg[0] (
	.clk(clk_clk),
	.d(\address_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[0]~q ),
	.prn(vcc));
defparam \address_reg[0] .is_wysiwyg = "true";
defparam \address_reg[0] .power_up = "low";

cycloneive_lcell_comb \readdata~1 (
	.dataa(\readdata~0_combout ),
	.datab(src_data_39),
	.datac(\address_reg[0]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hFEFF;
defparam \readdata~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~2 (
	.dataa(readdata_0),
	.datab(\readdata~1_combout ),
	.datac(gnd),
	.datad(m0_read),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hAACC;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg~3 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_reg~3_combout ),
	.cout());
defparam \control_reg~3 .lut_mask = 16'hFBFB;
defparam \control_reg~3 .sum_lutc_input = "datac";

dffeas \address_reg[1] (
	.clk(clk_clk),
	.d(\control_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[1]~q ),
	.prn(vcc));
defparam \address_reg[1] .is_wysiwyg = "true";
defparam \address_reg[1] .power_up = "low";

cycloneive_lcell_comb \internal_reset~3 (
	.dataa(d_writedata_0),
	.datab(src_data_32),
	.datac(src_data_38),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\internal_reset~3_combout ),
	.cout());
defparam \internal_reset~3 .lut_mask = 16'hEFFF;
defparam \internal_reset~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~12 (
	.dataa(internal_reset),
	.datab(\internal_reset~3_combout ),
	.datac(r_sync_rst),
	.datad(\Serial_Bus_Controller|transfer_complete~q ),
	.cin(gnd),
	.combout(\s_serial_transfer~12_combout ),
	.cout());
defparam \s_serial_transfer~12 .lut_mask = 16'h7FFF;
defparam \s_serial_transfer~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\s_serial_transfer.STATE_4_PRE_READ~q ),
	.datab(\s_serial_transfer.STATE_5_READ_TRANSFER~q ),
	.datac(gnd),
	.datad(\Serial_Bus_Controller|transfer_complete~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_5_READ_TRANSFER (
	.clk(clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_transfer.STATE_5_READ_TRANSFER~q ),
	.prn(vcc));
defparam \s_serial_transfer.STATE_5_READ_TRANSFER .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_5_READ_TRANSFER .power_up = "low";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\Serial_Bus_Controller|transfer_complete~q ),
	.datab(\s_serial_transfer.STATE_5_READ_TRANSFER~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hEEEE;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg[17]~0 (
	.dataa(s_serial_transferSTATE_1_PRE_WRITE),
	.datab(Equal2),
	.datac(saved_grant_1),
	.datad(d_byteenable_2),
	.cin(gnd),
	.combout(\control_reg[17]~0_combout ),
	.cout());
defparam \control_reg[17]~0 .lut_mask = 16'hDFFF;
defparam \control_reg[17]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg[17]~1 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(\control_reg[17]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_reg[17]~1_combout ),
	.cout());
defparam \control_reg[17]~1 .lut_mask = 16'hFEFE;
defparam \control_reg[17]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg[17]~2 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(internal_reset),
	.datac(waitrequest1),
	.datad(\control_reg[17]~1_combout ),
	.cin(gnd),
	.combout(\control_reg[17]~2_combout ),
	.cout());
defparam \control_reg[17]~2 .lut_mask = 16'hEFFF;
defparam \control_reg[17]~2 .sum_lutc_input = "datac";

dffeas \control_reg[16] (
	.clk(clk_clk),
	.d(src_payload),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(\control_reg[17]~2_combout ),
	.q(\control_reg[16]~q ),
	.prn(vcc));
defparam \control_reg[16] .is_wysiwyg = "true";
defparam \control_reg[16] .power_up = "low";

dffeas \control_reg[17] (
	.clk(clk_clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(\control_reg[17]~2_combout ),
	.q(\control_reg[17]~q ),
	.prn(vcc));
defparam \control_reg[17] .is_wysiwyg = "true";
defparam \control_reg[17] .power_up = "low";

cycloneive_lcell_comb \Selector3~1 (
	.dataa(\Selector3~0_combout ),
	.datab(\s_serial_transfer~14_combout ),
	.datac(\control_reg[16]~q ),
	.datad(\control_reg[17]~q ),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'hEFFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_6_POST_READ (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_transfer.STATE_6_POST_READ~q ),
	.prn(vcc));
defparam \s_serial_transfer.STATE_6_POST_READ .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_6_POST_READ .power_up = "low";

cycloneive_lcell_comb \ns_serial_transfer~2 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(\AV_Config_Auto_Init|auto_init_complete~q ),
	.datad(\Serial_Bus_Controller|transfer_complete~q ),
	.cin(gnd),
	.combout(\ns_serial_transfer~2_combout ),
	.cout());
defparam \ns_serial_transfer~2 .lut_mask = 16'hFEFF;
defparam \ns_serial_transfer~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~18 (
	.dataa(saved_grant_0),
	.datab(uav_write),
	.datac(src_data_68),
	.datad(\ns_serial_transfer~2_combout ),
	.cin(gnd),
	.combout(\s_serial_transfer~18_combout ),
	.cout());
defparam \s_serial_transfer~18 .lut_mask = 16'h7FFF;
defparam \s_serial_transfer~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~19 (
	.dataa(mem_used_1),
	.datab(\s_serial_transfer~18_combout ),
	.datac(WideOr1),
	.datad(\s_serial_transfer.STATE_0_IDLE~q ),
	.cin(gnd),
	.combout(\s_serial_transfer~19_combout ),
	.cout());
defparam \s_serial_transfer~19 .lut_mask = 16'hEFFF;
defparam \s_serial_transfer~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(s_serial_transferSTATE_1_PRE_WRITE),
	.datab(\s_serial_transfer.STATE_2_WRITE_TRANSFER~q ),
	.datac(gnd),
	.datad(\Serial_Bus_Controller|transfer_complete~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hEEFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_2_WRITE_TRANSFER (
	.clk(clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_transfer.STATE_2_WRITE_TRANSFER~q ),
	.prn(vcc));
defparam \s_serial_transfer.STATE_2_WRITE_TRANSFER .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_2_WRITE_TRANSFER .power_up = "low";

cycloneive_lcell_comb \s_serial_transfer~21 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(\Serial_Bus_Controller|transfer_complete~q ),
	.datac(\s_serial_transfer.STATE_2_WRITE_TRANSFER~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\s_serial_transfer~21_combout ),
	.cout());
defparam \s_serial_transfer~21 .lut_mask = 16'hFDFD;
defparam \s_serial_transfer~21 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_3_POST_WRITE (
	.clk(clk_clk),
	.d(\s_serial_transfer~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_transfer.STATE_3_POST_WRITE~q ),
	.prn(vcc));
defparam \s_serial_transfer.STATE_3_POST_WRITE .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_3_POST_WRITE .power_up = "low";

cycloneive_lcell_comb \s_serial_transfer~20 (
	.dataa(\s_serial_transfer.STATE_6_POST_READ~q ),
	.datab(\s_serial_transfer~19_combout ),
	.datac(\s_serial_transfer.STATE_3_POST_WRITE~q ),
	.datad(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.cin(gnd),
	.combout(\s_serial_transfer~20_combout ),
	.cout());
defparam \s_serial_transfer~20 .lut_mask = 16'h7FFF;
defparam \s_serial_transfer~20 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_0_IDLE (
	.clk(clk_clk),
	.d(\s_serial_transfer~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_transfer.STATE_0_IDLE~q ),
	.prn(vcc));
defparam \s_serial_transfer.STATE_0_IDLE .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_0_IDLE .power_up = "low";

cycloneive_lcell_comb \s_serial_transfer~13 (
	.dataa(\AV_Config_Auto_Init|auto_init_complete~q ),
	.datab(Equal2),
	.datac(\Serial_Bus_Controller|transfer_complete~q ),
	.datad(\s_serial_transfer.STATE_0_IDLE~q ),
	.cin(gnd),
	.combout(\s_serial_transfer~13_combout ),
	.cout());
defparam \s_serial_transfer~13 .lut_mask = 16'hEFFF;
defparam \s_serial_transfer~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~14 (
	.dataa(\s_serial_transfer~13_combout ),
	.datab(internal_reset),
	.datac(Equal2),
	.datad(m0_read),
	.cin(gnd),
	.combout(\s_serial_transfer~14_combout ),
	.cout());
defparam \s_serial_transfer~14 .lut_mask = 16'hBFFF;
defparam \s_serial_transfer~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~17 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(\s_serial_transfer~14_combout ),
	.datac(\control_reg[16]~q ),
	.datad(\control_reg[17]~q ),
	.cin(gnd),
	.combout(\s_serial_transfer~17_combout ),
	.cout());
defparam \s_serial_transfer~17 .lut_mask = 16'hFFFD;
defparam \s_serial_transfer~17 .sum_lutc_input = "datac";

dffeas \s_serial_transfer.STATE_4_PRE_READ (
	.clk(clk_clk),
	.d(\s_serial_transfer~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_transfer.STATE_4_PRE_READ~q ),
	.prn(vcc));
defparam \s_serial_transfer.STATE_4_PRE_READ .is_wysiwyg = "true";
defparam \s_serial_transfer.STATE_4_PRE_READ .power_up = "low";

cycloneive_lcell_comb \start_external_transfer~0 (
	.dataa(s_serial_transferSTATE_1_PRE_WRITE),
	.datab(\s_serial_transfer.STATE_4_PRE_READ~q ),
	.datac(gnd),
	.datad(\s_serial_transfer~12_combout ),
	.cin(gnd),
	.combout(\start_external_transfer~0_combout ),
	.cout());
defparam \start_external_transfer~0 .lut_mask = 16'hEEFF;
defparam \start_external_transfer~0 .sum_lutc_input = "datac";

dffeas start_external_transfer(
	.clk(clk_clk),
	.d(\s_serial_transfer~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\start_external_transfer~0_combout ),
	.q(\start_external_transfer~q ),
	.prn(vcc));
defparam start_external_transfer.is_wysiwyg = "true";
defparam start_external_transfer.power_up = "low";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\AV_Config_Auto_Init|auto_init_complete~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\start_external_transfer~q ),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hAAFF;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg[2]~4 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(src_data_32),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_reg[2]~4_combout ),
	.cout());
defparam \control_reg[2]~4 .lut_mask = 16'hEFEF;
defparam \control_reg[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg[2]~5 (
	.dataa(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datab(internal_reset),
	.datac(waitrequest2),
	.datad(\control_reg[2]~4_combout ),
	.cin(gnd),
	.combout(\control_reg[2]~5_combout ),
	.cout());
defparam \control_reg[2]~5 .lut_mask = 16'hEFFF;
defparam \control_reg[2]~5 .sum_lutc_input = "datac";

dffeas \control_reg[1] (
	.clk(clk_clk),
	.d(\control_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_reg[2]~5_combout ),
	.q(\control_reg[1]~q ),
	.prn(vcc));
defparam \control_reg[1] .is_wysiwyg = "true";
defparam \control_reg[1] .power_up = "low";

cycloneive_lcell_comb \readdata~4 (
	.dataa(src_data_39),
	.datab(\readdata~3_combout ),
	.datac(src_data_38),
	.datad(\control_reg[1]~q ),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hFFDE;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\address_reg[1]~q ),
	.datab(src_data_39),
	.datac(\readdata~4_combout ),
	.datad(\Serial_Bus_Controller|shiftreg_data[2]~q ),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hFFBE;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(readdata_1),
	.datab(\readdata~5_combout ),
	.datac(gnd),
	.datad(m0_read),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hAACC;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(\Serial_Bus_Controller|shiftreg_data[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hFEFE;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \control_reg~6 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_reg~6_combout ),
	.cout());
defparam \control_reg~6 .lut_mask = 16'hFBFB;
defparam \control_reg~6 .sum_lutc_input = "datac";

dffeas \address_reg[2] (
	.clk(clk_clk),
	.d(\control_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[2]~q ),
	.prn(vcc));
defparam \address_reg[2] .is_wysiwyg = "true";
defparam \address_reg[2] .power_up = "low";

dffeas \control_reg[2] (
	.clk(clk_clk),
	.d(\control_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_reg[2]~5_combout ),
	.q(\control_reg[2]~q ),
	.prn(vcc));
defparam \control_reg[2] .is_wysiwyg = "true";
defparam \control_reg[2] .power_up = "low";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\address_reg[2]~q ),
	.datab(\control_reg[2]~q ),
	.datac(src_data_39),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hACFF;
defparam \readdata~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~9 (
	.dataa(readdata_2),
	.datab(\readdata~7_combout ),
	.datac(\readdata~8_combout ),
	.datad(m0_read),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hFAFC;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(src_data_38),
	.datab(\control_reg[16]~q ),
	.datac(gnd),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hEEFF;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3]~12 (
	.dataa(m0_read),
	.datab(internal_reset),
	.datac(\internal_reset~3_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[3]~12_combout ),
	.cout());
defparam \readdata[3]~12 .lut_mask = 16'hFFFD;
defparam \readdata[3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(src_data_38),
	.datab(\control_reg[17]~q ),
	.datac(gnd),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hEEFF;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\Serial_Bus_Controller|shiftreg_data[10]~q ),
	.datab(gnd),
	.datac(\control_reg[16]~q ),
	.datad(\control_reg[17]~q ),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hAFFF;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(\readdata~17_combout ),
	.datab(src_data_39),
	.datac(\AV_Config_Auto_Init|auto_init_complete~q ),
	.datad(\AV_Config_Auto_Init|auto_init_error~q ),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hB8FF;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(readdata_8),
	.datab(src_data_38),
	.datac(\readdata~18_combout ),
	.datad(m0_read),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hFAFC;
defparam \readdata~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_reset~4 (
	.dataa(d_write),
	.datab(write_accepted),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\internal_reset~4_combout ),
	.cout());
defparam \internal_reset~4 .lut_mask = 16'hFBFF;
defparam \internal_reset~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \waitrequest~0 (
	.dataa(src_data_38),
	.datab(src_data_39),
	.datac(gnd),
	.datad(\s_serial_transfer.STATE_6_POST_READ~q ),
	.cin(gnd),
	.combout(\waitrequest~0_combout ),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hEEFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~15 (
	.dataa(\AV_Config_Auto_Init|auto_init_complete~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\s_serial_transfer.STATE_0_IDLE~q ),
	.cin(gnd),
	.combout(\s_serial_transfer~15_combout ),
	.cout());
defparam \s_serial_transfer~15 .lut_mask = 16'hAAFF;
defparam \s_serial_transfer~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_transfer~16 (
	.dataa(internal_reset),
	.datab(Equal2),
	.datac(\s_serial_transfer~12_combout ),
	.datad(\s_serial_transfer~15_combout ),
	.cin(gnd),
	.combout(\s_serial_transfer~16_combout ),
	.cout());
defparam \s_serial_transfer~16 .lut_mask = 16'hFFFE;
defparam \s_serial_transfer~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3]~10 (
	.dataa(src_data_39),
	.datab(internal_reset),
	.datac(\internal_reset~3_combout ),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\readdata[3]~10_combout ),
	.cout());
defparam \readdata[3]~10 .lut_mask = 16'hBFFF;
defparam \readdata[3]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~3 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg~3_combout ),
	.cout());
defparam \address_reg~3 .lut_mask = 16'hFBFB;
defparam \address_reg~3 .sum_lutc_input = "datac";

dffeas \address_reg[3] (
	.clk(clk_clk),
	.d(\address_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[3]~q ),
	.prn(vcc));
defparam \address_reg[3] .is_wysiwyg = "true";
defparam \address_reg[3] .power_up = "low";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\readdata[3]~10_combout ),
	.datab(\Serial_Bus_Controller|shiftreg_data[4]~q ),
	.datac(\address_reg[3]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hFAFC;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~4 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg~4_combout ),
	.cout());
defparam \address_reg~4 .lut_mask = 16'hFBFB;
defparam \address_reg~4 .sum_lutc_input = "datac";

dffeas \address_reg[4] (
	.clk(clk_clk),
	.d(\address_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[4]~q ),
	.prn(vcc));
defparam \address_reg[4] .is_wysiwyg = "true";
defparam \address_reg[4] .power_up = "low";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\readdata[3]~10_combout ),
	.datab(\Serial_Bus_Controller|shiftreg_data[5]~q ),
	.datac(\address_reg[4]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hFAFC;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~5 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg~5_combout ),
	.cout());
defparam \address_reg~5 .lut_mask = 16'hFBFB;
defparam \address_reg~5 .sum_lutc_input = "datac";

dffeas \address_reg[5] (
	.clk(clk_clk),
	.d(\address_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[5]~q ),
	.prn(vcc));
defparam \address_reg[5] .is_wysiwyg = "true";
defparam \address_reg[5] .power_up = "low";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\readdata[3]~10_combout ),
	.datab(\Serial_Bus_Controller|shiftreg_data[6]~q ),
	.datac(\address_reg[5]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hFAFC;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~6 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg~6_combout ),
	.cout());
defparam \address_reg~6 .lut_mask = 16'hFBFB;
defparam \address_reg~6 .sum_lutc_input = "datac";

dffeas \address_reg[7] (
	.clk(clk_clk),
	.d(\address_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[7]~q ),
	.prn(vcc));
defparam \address_reg[7] .is_wysiwyg = "true";
defparam \address_reg[7] .power_up = "low";

cycloneive_lcell_comb \readdata~20 (
	.dataa(\readdata[3]~10_combout ),
	.datab(\Serial_Bus_Controller|shiftreg_data[8]~q ),
	.datac(\address_reg[7]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hFAFC;
defparam \readdata~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \address_reg~7 (
	.dataa(saved_grant_0),
	.datab(\Serial_Bus_Controller|shiftreg_mask~2_combout ),
	.datac(d_writedata_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg~7_combout ),
	.cout());
defparam \address_reg~7 .lut_mask = 16'hFBFB;
defparam \address_reg~7 .sum_lutc_input = "datac";

dffeas \address_reg[6] (
	.clk(clk_clk),
	.d(\address_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg[4]~2_combout ),
	.q(\address_reg[6]~q ),
	.prn(vcc));
defparam \address_reg[6] .is_wysiwyg = "true";
defparam \address_reg[6] .power_up = "low";

cycloneive_lcell_comb \readdata~21 (
	.dataa(\readdata[3]~10_combout ),
	.datab(\Serial_Bus_Controller|shiftreg_data[7]~q ),
	.datac(\address_reg[6]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hFAFC;
defparam \readdata~21 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_av_config_auto_init (
	transfer_data1,
	auto_init_complete1,
	transfer_complete,
	rom_address_4,
	rom_address_1,
	rom_address_0,
	rom_address_2,
	rom_address_3,
	rom_address_5,
	data_out_25,
	auto_init_error1,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_10,
	data_out_8,
	data_out_7,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_out_12,
	data_out_11,
	shiftreg_mask,
	Ram0,
	ack,
	Ram01,
	data_out_24,
	rom_data_2,
	rom_data_3,
	rom_data_4,
	rom_data_5,
	WideOr0,
	rom_data_6,
	Ram02,
	rom_data_8,
	rom_data_7,
	Ram03,
	Ram04,
	Ram05,
	rom_data_14,
	rom_data_13,
	rom_data_11,
	rom_data_1,
	rom_data_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	transfer_data1;
output 	auto_init_complete1;
input 	transfer_complete;
output 	rom_address_4;
output 	rom_address_1;
output 	rom_address_0;
output 	rom_address_2;
output 	rom_address_3;
output 	rom_address_5;
output 	data_out_25;
output 	auto_init_error1;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_10;
output 	data_out_8;
output 	data_out_7;
output 	data_out_17;
output 	data_out_16;
output 	data_out_15;
output 	data_out_14;
output 	data_out_13;
output 	data_out_12;
output 	data_out_11;
input 	shiftreg_mask;
input 	Ram0;
input 	ack;
input 	Ram01;
output 	data_out_24;
input 	rom_data_2;
input 	rom_data_3;
input 	rom_data_4;
input 	rom_data_5;
input 	WideOr0;
input 	rom_data_6;
input 	Ram02;
input 	rom_data_8;
input 	rom_data_7;
input 	Ram03;
input 	Ram04;
input 	Ram05;
input 	rom_data_14;
input 	rom_data_13;
input 	rom_data_11;
input 	rom_data_1;
input 	rom_data_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always1~0_combout ;
wire \always3~0_combout ;
wire \auto_init_complete~0_combout ;
wire \rom_address[0]~7 ;
wire \rom_address[1]~9 ;
wire \rom_address[2]~11 ;
wire \rom_address[3]~13 ;
wire \rom_address[4]~14_combout ;
wire \rom_address[4]~16_combout ;
wire \rom_address[1]~8_combout ;
wire \rom_address[0]~6_combout ;
wire \rom_address[2]~10_combout ;
wire \rom_address[3]~12_combout ;
wire \rom_address[4]~15 ;
wire \rom_address[5]~17_combout ;
wire \auto_init_error~0_combout ;
wire \data_out~0_combout ;


dffeas transfer_data(
	.clk(clk_clk),
	.d(\always1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(transfer_data1),
	.prn(vcc));
defparam transfer_data.is_wysiwyg = "true";
defparam transfer_data.power_up = "low";

dffeas auto_init_complete(
	.clk(clk_clk),
	.d(\auto_init_complete~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(auto_init_complete1),
	.prn(vcc));
defparam auto_init_complete.is_wysiwyg = "true";
defparam auto_init_complete.power_up = "low";

dffeas \rom_address[4] (
	.clk(clk_clk),
	.d(\rom_address[4]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\rom_address[4]~16_combout ),
	.q(rom_address_4),
	.prn(vcc));
defparam \rom_address[4] .is_wysiwyg = "true";
defparam \rom_address[4] .power_up = "low";

dffeas \rom_address[1] (
	.clk(clk_clk),
	.d(\rom_address[1]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\rom_address[4]~16_combout ),
	.q(rom_address_1),
	.prn(vcc));
defparam \rom_address[1] .is_wysiwyg = "true";
defparam \rom_address[1] .power_up = "low";

dffeas \rom_address[0] (
	.clk(clk_clk),
	.d(\rom_address[0]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\rom_address[4]~16_combout ),
	.q(rom_address_0),
	.prn(vcc));
defparam \rom_address[0] .is_wysiwyg = "true";
defparam \rom_address[0] .power_up = "low";

dffeas \rom_address[2] (
	.clk(clk_clk),
	.d(\rom_address[2]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\rom_address[4]~16_combout ),
	.q(rom_address_2),
	.prn(vcc));
defparam \rom_address[2] .is_wysiwyg = "true";
defparam \rom_address[2] .power_up = "low";

dffeas \rom_address[3] (
	.clk(clk_clk),
	.d(\rom_address[3]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\rom_address[4]~16_combout ),
	.q(rom_address_3),
	.prn(vcc));
defparam \rom_address[3] .is_wysiwyg = "true";
defparam \rom_address[3] .power_up = "low";

dffeas \rom_address[5] (
	.clk(clk_clk),
	.d(\rom_address[5]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\rom_address[4]~16_combout ),
	.q(rom_address_5),
	.prn(vcc));
defparam \rom_address[5] .is_wysiwyg = "true";
defparam \rom_address[5] .power_up = "low";

dffeas \data_out[25] (
	.clk(clk_clk),
	.d(Ram01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_25),
	.prn(vcc));
defparam \data_out[25] .is_wysiwyg = "true";
defparam \data_out[25] .power_up = "low";

dffeas auto_init_error(
	.clk(clk_clk),
	.d(\auto_init_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(auto_init_error1),
	.prn(vcc));
defparam auto_init_error.is_wysiwyg = "true";
defparam auto_init_error.power_up = "low";

dffeas \data_out[1] (
	.clk(clk_clk),
	.d(rom_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk_clk),
	.d(rom_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk_clk),
	.d(rom_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk_clk),
	.d(rom_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk_clk),
	.d(rom_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk_clk),
	.d(rom_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk_clk),
	.d(Ram02),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk_clk),
	.d(rom_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk_clk),
	.d(rom_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk_clk),
	.d(Ram03),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk_clk),
	.d(Ram04),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk_clk),
	.d(Ram05),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk_clk),
	.d(rom_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk_clk),
	.d(rom_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk_clk),
	.d(rom_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk_clk),
	.d(rom_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[24] (
	.clk(clk_clk),
	.d(\data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_24),
	.prn(vcc));
defparam \data_out[24] .is_wysiwyg = "true";
defparam \data_out[24] .power_up = "low";

cycloneive_lcell_comb \always1~0 (
	.dataa(transfer_complete),
	.datab(auto_init_complete1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'h7777;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always3~0 (
	.dataa(transfer_complete),
	.datab(transfer_data1),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hFFFE;
defparam \always3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_init_complete~0 (
	.dataa(auto_init_complete1),
	.datab(Ram0),
	.datac(\always3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_init_complete~0_combout ),
	.cout());
defparam \auto_init_complete~0 .lut_mask = 16'hFEFE;
defparam \auto_init_complete~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_address[0]~6 (
	.dataa(rom_address_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\rom_address[0]~6_combout ),
	.cout(\rom_address[0]~7 ));
defparam \rom_address[0]~6 .lut_mask = 16'h55AA;
defparam \rom_address[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_address[1]~8 (
	.dataa(rom_address_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rom_address[0]~7 ),
	.combout(\rom_address[1]~8_combout ),
	.cout(\rom_address[1]~9 ));
defparam \rom_address[1]~8 .lut_mask = 16'h5A5F;
defparam \rom_address[1]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \rom_address[2]~10 (
	.dataa(rom_address_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rom_address[1]~9 ),
	.combout(\rom_address[2]~10_combout ),
	.cout(\rom_address[2]~11 ));
defparam \rom_address[2]~10 .lut_mask = 16'h5AAF;
defparam \rom_address[2]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \rom_address[3]~12 (
	.dataa(rom_address_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rom_address[2]~11 ),
	.combout(\rom_address[3]~12_combout ),
	.cout(\rom_address[3]~13 ));
defparam \rom_address[3]~12 .lut_mask = 16'h5A5F;
defparam \rom_address[3]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \rom_address[4]~14 (
	.dataa(rom_address_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rom_address[3]~13 ),
	.combout(\rom_address[4]~14_combout ),
	.cout(\rom_address[4]~15 ));
defparam \rom_address[4]~14 .lut_mask = 16'h5AAF;
defparam \rom_address[4]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \rom_address[4]~16 (
	.dataa(shiftreg_mask),
	.datab(gnd),
	.datac(transfer_complete),
	.datad(transfer_data1),
	.cin(gnd),
	.combout(\rom_address[4]~16_combout ),
	.cout());
defparam \rom_address[4]~16 .lut_mask = 16'hFFFA;
defparam \rom_address[4]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_address[5]~17 (
	.dataa(rom_address_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\rom_address[4]~15 ),
	.combout(\rom_address[5]~17_combout ),
	.cout());
defparam \rom_address[5]~17 .lut_mask = 16'h5A5A;
defparam \rom_address[5]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_init_error~0 (
	.dataa(auto_init_error1),
	.datab(transfer_complete),
	.datac(transfer_data1),
	.datad(ack),
	.cin(gnd),
	.combout(\auto_init_error~0_combout ),
	.cout());
defparam \auto_init_error~0 .lut_mask = 16'hFFFE;
defparam \auto_init_error~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out~0 (
	.dataa(rom_address_5),
	.datab(WideOr0),
	.datac(gnd),
	.datad(shiftreg_mask),
	.cin(gnd),
	.combout(\data_out~0_combout ),
	.cout());
defparam \data_out~0 .lut_mask = 16'h77FF;
defparam \data_out~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_av_config_auto_init_ob_de2_115 (
	rom_address_4,
	rom_address_1,
	rom_address_0,
	rom_address_2,
	rom_address_3,
	rom_address_5,
	Ram0,
	Ram01,
	rom_data_2,
	rom_data_3,
	rom_data_4,
	rom_data_5,
	WideOr0,
	rom_data_6,
	Ram02,
	rom_data_8,
	rom_data_7,
	Ram03,
	Ram04,
	Ram05,
	rom_data_14,
	rom_data_13,
	rom_data_11,
	rom_data_1,
	rom_data_12)/* synthesis synthesis_greybox=1 */;
input 	rom_address_4;
input 	rom_address_1;
input 	rom_address_0;
input 	rom_address_2;
input 	rom_address_3;
input 	rom_address_5;
output 	Ram0;
output 	Ram01;
output 	rom_data_2;
output 	rom_data_3;
output 	rom_data_4;
output 	rom_data_5;
output 	WideOr0;
output 	rom_data_6;
output 	Ram02;
output 	rom_data_8;
output 	rom_data_7;
output 	Ram03;
output 	Ram04;
output 	Ram05;
output 	rom_data_14;
output 	rom_data_13;
output 	rom_data_11;
output 	rom_data_1;
output 	rom_data_12;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Auto_Init_Audio_ROM|Decoder0~0_combout ;
wire \Auto_Init_Audio_ROM|Decoder0~1_combout ;
wire \Auto_Init_Audio_ROM|Decoder0~2_combout ;
wire \Auto_Init_Video_ROM|Ram0~8_combout ;
wire \Auto_Init_Audio_ROM|Decoder0~3_combout ;
wire \Auto_Init_Video_ROM|Ram0~9_combout ;
wire \Auto_Init_Video_ROM|Ram0~16_combout ;
wire \Auto_Init_Video_ROM|Ram0~17_combout ;
wire \Auto_Init_Video_ROM|Ram0~18_combout ;
wire \rom_data[2]~38_combout ;
wire \rom_data[2]~39_combout ;
wire \rom_data[2]~40_combout ;
wire \rom_data[2]~41_combout ;
wire \rom_data[2]~42_combout ;
wire \rom_data[2]~43_combout ;
wire \rom_data[2]~44_combout ;
wire \rom_data[3]~46_combout ;
wire \rom_data[3]~47_combout ;
wire \rom_data[3]~48_combout ;
wire \rom_data[3]~49_combout ;
wire \rom_data[3]~50_combout ;
wire \rom_data[3]~51_combout ;
wire \rom_data[5]~53_combout ;
wire \rom_data[5]~54_combout ;
wire \rom_data[5]~55_combout ;
wire \rom_data[5]~56_combout ;
wire \rom_data[6]~3_combout ;
wire \rom_data[6]~4_combout ;
wire \rom_data[6]~78_combout ;
wire \rom_data[8]~59_combout ;
wire \rom_data[8]~60_combout ;
wire \rom_data[7]~37_combout ;
wire \rom_data[7]~62_combout ;
wire \rom_data[7]~63_combout ;
wire \rom_data[7]~64_combout ;
wire \rom_data[7]~65_combout ;
wire \rom_data[7]~66_combout ;
wire \rom_data[14]~68_combout ;
wire \rom_data[14]~69_combout ;
wire \rom_data[14]~70_combout ;
wire \rom_data[14]~71_combout ;
wire \rom_data[13]~73_combout ;
wire \rom_data[13]~74_combout ;
wire \rom_data[13]~75_combout ;
wire \rom_data[13]~76_combout ;
wire \rom_data[11]~13_combout ;
wire \rom_data[11]~11_combout ;
wire \rom_data[11]~10_combout ;
wire \rom_data[11]~31_combout ;
wire \rom_data[11]~14_combout ;
wire \rom_data[1]~21_combout ;
wire \rom_data[1]~19_combout ;
wire \rom_data[1]~18_combout ;
wire \rom_data[1]~33_combout ;
wire \rom_data[1]~22_combout ;
wire \rom_data[12]~29_combout ;
wire \rom_data[12]~27_combout ;
wire \rom_data[12]~26_combout ;
wire \rom_data[12]~35_combout ;
wire \rom_data[12]~30_combout ;


final_project_soc_altera_up_av_config_auto_init_ob_adv7180 Auto_Init_Video_ROM(
	.rom_address_4(rom_address_4),
	.rom_address_1(rom_address_1),
	.rom_address_0(rom_address_0),
	.rom_address_2(rom_address_2),
	.rom_address_3(rom_address_3),
	.rom_address_5(rom_address_5),
	.Ram0(Ram0),
	.Ram01(Ram01),
	.Ram02(\Auto_Init_Video_ROM|Ram0~8_combout ),
	.Ram03(\Auto_Init_Video_ROM|Ram0~9_combout ),
	.Ram04(Ram02),
	.Ram05(\Auto_Init_Video_ROM|Ram0~16_combout ),
	.Ram06(\Auto_Init_Video_ROM|Ram0~17_combout ),
	.Ram07(\Auto_Init_Video_ROM|Ram0~18_combout ),
	.Ram08(Ram03),
	.Ram09(Ram04),
	.Ram010(Ram05));

final_project_soc_altera_up_av_config_auto_init_ob_audio Auto_Init_Audio_ROM(
	.rom_address_4(rom_address_4),
	.rom_address_1(rom_address_1),
	.rom_address_0(rom_address_0),
	.rom_address_2(rom_address_2),
	.rom_address_3(rom_address_3),
	.rom_address_5(rom_address_5),
	.Decoder0(\Auto_Init_Audio_ROM|Decoder0~0_combout ),
	.Decoder01(\Auto_Init_Audio_ROM|Decoder0~1_combout ),
	.Decoder02(\Auto_Init_Audio_ROM|Decoder0~2_combout ),
	.Decoder03(\Auto_Init_Audio_ROM|Decoder0~3_combout ),
	.WideOr0(WideOr0));

cycloneive_lcell_comb \rom_data[2]~45 (
	.dataa(\rom_data[2]~38_combout ),
	.datab(\rom_data[2]~39_combout ),
	.datac(\rom_data[2]~43_combout ),
	.datad(\rom_data[2]~44_combout ),
	.cin(gnd),
	.combout(rom_data_2),
	.cout());
defparam \rom_data[2]~45 .lut_mask = 16'hF7D5;
defparam \rom_data[2]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~52 (
	.dataa(\rom_data[3]~46_combout ),
	.datab(\rom_data[3]~47_combout ),
	.datac(\rom_data[3]~50_combout ),
	.datad(\rom_data[3]~51_combout ),
	.cin(gnd),
	.combout(rom_data_3),
	.cout());
defparam \rom_data[3]~52 .lut_mask = 16'hF7D5;
defparam \rom_data[3]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[4] (
	.dataa(\Auto_Init_Video_ROM|Ram0~8_combout ),
	.datab(\Auto_Init_Audio_ROM|Decoder0~0_combout ),
	.datac(\Auto_Init_Audio_ROM|Decoder0~3_combout ),
	.datad(\rom_data[2]~38_combout ),
	.cin(gnd),
	.combout(rom_data_4),
	.cout());
defparam \rom_data[4] .lut_mask = 16'hFEFF;
defparam \rom_data[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[5]~57 (
	.dataa(\rom_data[2]~38_combout ),
	.datab(\rom_data[5]~53_combout ),
	.datac(\rom_data[5]~55_combout ),
	.datad(\rom_data[5]~56_combout ),
	.cin(gnd),
	.combout(rom_data_5),
	.cout());
defparam \rom_data[5]~57 .lut_mask = 16'hF7D5;
defparam \rom_data[5]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[6]~58 (
	.dataa(\rom_data[6]~78_combout ),
	.datab(rom_address_4),
	.datac(\Auto_Init_Video_ROM|Ram0~9_combout ),
	.datad(rom_address_1),
	.cin(gnd),
	.combout(rom_data_6),
	.cout());
defparam \rom_data[6]~58 .lut_mask = 16'hFEFF;
defparam \rom_data[6]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[8]~61 (
	.dataa(\rom_data[8]~60_combout ),
	.datab(\Auto_Init_Audio_ROM|Decoder0~2_combout ),
	.datac(rom_address_1),
	.datad(rom_address_0),
	.cin(gnd),
	.combout(rom_data_8),
	.cout());
defparam \rom_data[8]~61 .lut_mask = 16'hEFFF;
defparam \rom_data[8]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~67 (
	.dataa(\rom_data[7]~37_combout ),
	.datab(\rom_data[7]~62_combout ),
	.datac(\rom_data[7]~65_combout ),
	.datad(\rom_data[7]~66_combout ),
	.cin(gnd),
	.combout(rom_data_7),
	.cout());
defparam \rom_data[7]~67 .lut_mask = 16'hD77D;
defparam \rom_data[7]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[14]~72 (
	.dataa(rom_address_4),
	.datab(\rom_data[14]~70_combout ),
	.datac(\rom_data[14]~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(rom_data_14),
	.cout());
defparam \rom_data[14]~72 .lut_mask = 16'h9696;
defparam \rom_data[14]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[13]~77 (
	.dataa(rom_address_3),
	.datab(\Auto_Init_Audio_ROM|Decoder0~2_combout ),
	.datac(\rom_data[13]~75_combout ),
	.datad(\rom_data[13]~76_combout ),
	.cin(gnd),
	.combout(rom_data_13),
	.cout());
defparam \rom_data[13]~77 .lut_mask = 16'hEDDE;
defparam \rom_data[13]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[11]~32 (
	.dataa(\rom_data[11]~13_combout ),
	.datab(rom_address_2),
	.datac(\rom_data[11]~31_combout ),
	.datad(\rom_data[11]~14_combout ),
	.cin(gnd),
	.combout(rom_data_11),
	.cout());
defparam \rom_data[11]~32 .lut_mask = 16'hFFBE;
defparam \rom_data[11]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[1]~34 (
	.dataa(\rom_data[1]~21_combout ),
	.datab(rom_address_2),
	.datac(\rom_data[1]~33_combout ),
	.datad(\rom_data[1]~22_combout ),
	.cin(gnd),
	.combout(rom_data_1),
	.cout());
defparam \rom_data[1]~34 .lut_mask = 16'hFFBE;
defparam \rom_data[1]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[12]~36 (
	.dataa(\rom_data[12]~29_combout ),
	.datab(rom_address_2),
	.datac(\rom_data[12]~35_combout ),
	.datad(\rom_data[12]~30_combout ),
	.cin(gnd),
	.combout(rom_data_12),
	.cout());
defparam \rom_data[12]~36 .lut_mask = 16'hFFBE;
defparam \rom_data[12]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~38 (
	.dataa(rom_address_2),
	.datab(rom_address_1),
	.datac(rom_address_0),
	.datad(\Auto_Init_Audio_ROM|Decoder0~1_combout ),
	.cin(gnd),
	.combout(\rom_data[2]~38_combout ),
	.cout());
defparam \rom_data[2]~38 .lut_mask = 16'hFEFF;
defparam \rom_data[2]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~39 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(rom_address_5),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[2]~39_combout ),
	.cout());
defparam \rom_data[2]~39 .lut_mask = 16'hFF96;
defparam \rom_data[2]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~40 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(rom_address_5),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[2]~40_combout ),
	.cout());
defparam \rom_data[2]~40 .lut_mask = 16'hD77D;
defparam \rom_data[2]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~41 (
	.dataa(rom_address_0),
	.datab(\Auto_Init_Audio_ROM|Decoder0~2_combout ),
	.datac(rom_address_1),
	.datad(\rom_data[2]~40_combout ),
	.cin(gnd),
	.combout(\rom_data[2]~41_combout ),
	.cout());
defparam \rom_data[2]~41 .lut_mask = 16'hFFDE;
defparam \rom_data[2]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~42 (
	.dataa(rom_address_0),
	.datab(\Auto_Init_Audio_ROM|Decoder0~2_combout ),
	.datac(rom_address_1),
	.datad(\rom_data[2]~40_combout ),
	.cin(gnd),
	.combout(\rom_data[2]~42_combout ),
	.cout());
defparam \rom_data[2]~42 .lut_mask = 16'hF7B3;
defparam \rom_data[2]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~43 (
	.dataa(rom_address_4),
	.datab(rom_address_0),
	.datac(\rom_data[2]~41_combout ),
	.datad(\rom_data[2]~42_combout ),
	.cin(gnd),
	.combout(\rom_data[2]~43_combout ),
	.cout());
defparam \rom_data[2]~43 .lut_mask = 16'h6996;
defparam \rom_data[2]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[2]~44 (
	.dataa(rom_address_4),
	.datab(rom_address_0),
	.datac(\rom_data[2]~41_combout ),
	.datad(\rom_data[2]~42_combout ),
	.cin(gnd),
	.combout(\rom_data[2]~44_combout ),
	.cout());
defparam \rom_data[2]~44 .lut_mask = 16'h6996;
defparam \rom_data[2]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~46 (
	.dataa(gnd),
	.datab(rom_address_0),
	.datac(rom_address_2),
	.datad(\Auto_Init_Audio_ROM|Decoder0~1_combout ),
	.cin(gnd),
	.combout(\rom_data[3]~46_combout ),
	.cout());
defparam \rom_data[3]~46 .lut_mask = 16'h3FFF;
defparam \rom_data[3]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~47 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[3]~47_combout ),
	.cout());
defparam \rom_data[3]~47 .lut_mask = 16'h6996;
defparam \rom_data[3]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~48 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[3]~48_combout ),
	.cout());
defparam \rom_data[3]~48 .lut_mask = 16'h6996;
defparam \rom_data[3]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~49 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[3]~49_combout ),
	.cout());
defparam \rom_data[3]~49 .lut_mask = 16'hFF96;
defparam \rom_data[3]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~50 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(\rom_data[3]~48_combout ),
	.datad(\rom_data[3]~49_combout ),
	.cin(gnd),
	.combout(\rom_data[3]~50_combout ),
	.cout());
defparam \rom_data[3]~50 .lut_mask = 16'h6996;
defparam \rom_data[3]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[3]~51 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(\rom_data[3]~48_combout ),
	.datad(\rom_data[3]~49_combout ),
	.cin(gnd),
	.combout(\rom_data[3]~51_combout ),
	.cout());
defparam \rom_data[3]~51 .lut_mask = 16'h6996;
defparam \rom_data[3]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[5]~53 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[5]~53_combout ),
	.cout());
defparam \rom_data[5]~53 .lut_mask = 16'hB77B;
defparam \rom_data[5]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[5]~54 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[5]~54_combout ),
	.cout());
defparam \rom_data[5]~54 .lut_mask = 16'h6996;
defparam \rom_data[5]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[5]~55 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_5),
	.datad(\rom_data[5]~54_combout ),
	.cin(gnd),
	.combout(\rom_data[5]~55_combout ),
	.cout());
defparam \rom_data[5]~55 .lut_mask = 16'h6996;
defparam \rom_data[5]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[5]~56 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_5),
	.datad(\rom_data[5]~54_combout ),
	.cin(gnd),
	.combout(\rom_data[5]~56_combout ),
	.cout());
defparam \rom_data[5]~56 .lut_mask = 16'h6996;
defparam \rom_data[5]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[6]~3 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[6]~3_combout ),
	.cout());
defparam \rom_data[6]~3 .lut_mask = 16'h6996;
defparam \rom_data[6]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[6]~4 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[6]~4_combout ),
	.cout());
defparam \rom_data[6]~4 .lut_mask = 16'h6996;
defparam \rom_data[6]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[6]~78 (
	.dataa(\rom_data[6]~3_combout ),
	.datab(\rom_data[6]~4_combout ),
	.datac(rom_address_4),
	.datad(rom_address_1),
	.cin(gnd),
	.combout(\rom_data[6]~78_combout ),
	.cout());
defparam \rom_data[6]~78 .lut_mask = 16'hFFAC;
defparam \rom_data[6]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[8]~59 (
	.dataa(rom_address_1),
	.datab(\Auto_Init_Video_ROM|Ram0~16_combout ),
	.datac(\Auto_Init_Video_ROM|Ram0~17_combout ),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\rom_data[8]~59_combout ),
	.cout());
defparam \rom_data[8]~59 .lut_mask = 16'hFAFC;
defparam \rom_data[8]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[8]~60 (
	.dataa(\rom_data[8]~59_combout ),
	.datab(rom_address_3),
	.datac(\Auto_Init_Video_ROM|Ram0~18_combout ),
	.datad(rom_address_1),
	.cin(gnd),
	.combout(\rom_data[8]~60_combout ),
	.cout());
defparam \rom_data[8]~60 .lut_mask = 16'hFEFF;
defparam \rom_data[8]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~37 (
	.dataa(rom_address_2),
	.datab(gnd),
	.datac(rom_address_0),
	.datad(\Auto_Init_Audio_ROM|Decoder0~0_combout ),
	.cin(gnd),
	.combout(\rom_data[7]~37_combout ),
	.cout());
defparam \rom_data[7]~37 .lut_mask = 16'hAFFF;
defparam \rom_data[7]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~62 (
	.dataa(rom_address_5),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_0),
	.cin(gnd),
	.combout(\rom_data[7]~62_combout ),
	.cout());
defparam \rom_data[7]~62 .lut_mask = 16'hF9F6;
defparam \rom_data[7]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~63 (
	.dataa(rom_address_5),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_0),
	.cin(gnd),
	.combout(\rom_data[7]~63_combout ),
	.cout());
defparam \rom_data[7]~63 .lut_mask = 16'hF9F6;
defparam \rom_data[7]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~64 (
	.dataa(rom_address_5),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_0),
	.cin(gnd),
	.combout(\rom_data[7]~64_combout ),
	.cout());
defparam \rom_data[7]~64 .lut_mask = 16'h6996;
defparam \rom_data[7]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~65 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(\rom_data[7]~63_combout ),
	.datad(\rom_data[7]~64_combout ),
	.cin(gnd),
	.combout(\rom_data[7]~65_combout ),
	.cout());
defparam \rom_data[7]~65 .lut_mask = 16'hEDDE;
defparam \rom_data[7]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[7]~66 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(\rom_data[7]~63_combout ),
	.datad(\rom_data[7]~64_combout ),
	.cin(gnd),
	.combout(\rom_data[7]~66_combout ),
	.cout());
defparam \rom_data[7]~66 .lut_mask = 16'hFFD8;
defparam \rom_data[7]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[14]~68 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[14]~68_combout ),
	.cout());
defparam \rom_data[14]~68 .lut_mask = 16'hFF96;
defparam \rom_data[14]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[14]~69 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[14]~69_combout ),
	.cout());
defparam \rom_data[14]~69 .lut_mask = 16'hF9F6;
defparam \rom_data[14]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[14]~70 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(\rom_data[14]~68_combout ),
	.datad(\rom_data[14]~69_combout ),
	.cin(gnd),
	.combout(\rom_data[14]~70_combout ),
	.cout());
defparam \rom_data[14]~70 .lut_mask = 16'h6996;
defparam \rom_data[14]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[14]~71 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(\rom_data[14]~68_combout ),
	.datad(\rom_data[14]~69_combout ),
	.cin(gnd),
	.combout(\rom_data[14]~71_combout ),
	.cout());
defparam \rom_data[14]~71 .lut_mask = 16'h6996;
defparam \rom_data[14]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[13]~73 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[13]~73_combout ),
	.cout());
defparam \rom_data[13]~73 .lut_mask = 16'hFFBE;
defparam \rom_data[13]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[13]~74 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[13]~74_combout ),
	.cout());
defparam \rom_data[13]~74 .lut_mask = 16'hFFFE;
defparam \rom_data[13]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[13]~75 (
	.dataa(rom_address_2),
	.datab(rom_address_4),
	.datac(\rom_data[13]~73_combout ),
	.datad(\rom_data[13]~74_combout ),
	.cin(gnd),
	.combout(\rom_data[13]~75_combout ),
	.cout());
defparam \rom_data[13]~75 .lut_mask = 16'hEDDE;
defparam \rom_data[13]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[13]~76 (
	.dataa(rom_address_2),
	.datab(rom_address_4),
	.datac(\rom_data[13]~73_combout ),
	.datad(\rom_data[13]~74_combout ),
	.cin(gnd),
	.combout(\rom_data[13]~76_combout ),
	.cout());
defparam \rom_data[13]~76 .lut_mask = 16'h6996;
defparam \rom_data[13]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[11]~13 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[11]~13_combout ),
	.cout());
defparam \rom_data[11]~13 .lut_mask = 16'h6996;
defparam \rom_data[11]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[11]~11 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[11]~11_combout ),
	.cout());
defparam \rom_data[11]~11 .lut_mask = 16'hF9F6;
defparam \rom_data[11]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[11]~10 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[11]~10_combout ),
	.cout());
defparam \rom_data[11]~10 .lut_mask = 16'h96FF;
defparam \rom_data[11]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[11]~31 (
	.dataa(rom_address_2),
	.datab(\rom_data[11]~11_combout ),
	.datac(rom_address_1),
	.datad(\rom_data[11]~10_combout ),
	.cin(gnd),
	.combout(\rom_data[11]~31_combout ),
	.cout());
defparam \rom_data[11]~31 .lut_mask = 16'hFFDE;
defparam \rom_data[11]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[11]~14 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[11]~14_combout ),
	.cout());
defparam \rom_data[11]~14 .lut_mask = 16'h6996;
defparam \rom_data[11]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[1]~21 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[1]~21_combout ),
	.cout());
defparam \rom_data[1]~21 .lut_mask = 16'h6996;
defparam \rom_data[1]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[1]~19 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[1]~19_combout ),
	.cout());
defparam \rom_data[1]~19 .lut_mask = 16'h6996;
defparam \rom_data[1]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[1]~18 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[1]~18_combout ),
	.cout());
defparam \rom_data[1]~18 .lut_mask = 16'h6996;
defparam \rom_data[1]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[1]~33 (
	.dataa(rom_address_2),
	.datab(\rom_data[1]~19_combout ),
	.datac(rom_address_1),
	.datad(\rom_data[1]~18_combout ),
	.cin(gnd),
	.combout(\rom_data[1]~33_combout ),
	.cout());
defparam \rom_data[1]~33 .lut_mask = 16'hFFDE;
defparam \rom_data[1]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[1]~22 (
	.dataa(rom_address_0),
	.datab(rom_address_3),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[1]~22_combout ),
	.cout());
defparam \rom_data[1]~22 .lut_mask = 16'h6996;
defparam \rom_data[1]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[12]~29 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[12]~29_combout ),
	.cout());
defparam \rom_data[12]~29 .lut_mask = 16'hDFEF;
defparam \rom_data[12]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[12]~27 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[12]~27_combout ),
	.cout());
defparam \rom_data[12]~27 .lut_mask = 16'hEFFF;
defparam \rom_data[12]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[12]~26 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[12]~26_combout ),
	.cout());
defparam \rom_data[12]~26 .lut_mask = 16'h6996;
defparam \rom_data[12]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[12]~35 (
	.dataa(rom_address_2),
	.datab(\rom_data[12]~27_combout ),
	.datac(rom_address_0),
	.datad(\rom_data[12]~26_combout ),
	.cin(gnd),
	.combout(\rom_data[12]~35_combout ),
	.cout());
defparam \rom_data[12]~35 .lut_mask = 16'hFFDE;
defparam \rom_data[12]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rom_data[12]~30 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\rom_data[12]~30_combout ),
	.cout());
defparam \rom_data[12]~30 .lut_mask = 16'h6996;
defparam \rom_data[12]~30 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_av_config_auto_init_ob_adv7180 (
	rom_address_4,
	rom_address_1,
	rom_address_0,
	rom_address_2,
	rom_address_3,
	rom_address_5,
	Ram0,
	Ram01,
	Ram02,
	Ram03,
	Ram04,
	Ram05,
	Ram06,
	Ram07,
	Ram08,
	Ram09,
	Ram010)/* synthesis synthesis_greybox=1 */;
input 	rom_address_4;
input 	rom_address_1;
input 	rom_address_0;
input 	rom_address_2;
input 	rom_address_3;
input 	rom_address_5;
output 	Ram0;
output 	Ram01;
output 	Ram02;
output 	Ram03;
output 	Ram04;
output 	Ram05;
output 	Ram06;
output 	Ram07;
output 	Ram08;
output 	Ram09;
output 	Ram010;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Ram0~1_combout ;
wire \Ram0~2_combout ;
wire \Ram0~4_combout ;
wire \Ram0~5_combout ;
wire \Ram0~6_combout ;
wire \Ram0~7_combout ;
wire \Ram0~10_combout ;
wire \Ram0~11_combout ;
wire \Ram0~12_combout ;
wire \Ram0~13_combout ;
wire \Ram0~14_combout ;
wire \Ram0~19_combout ;
wire \Ram0~21_combout ;
wire \Ram0~23_combout ;
wire \Ram0~24_combout ;


cycloneive_lcell_comb \Ram0~0 (
	.dataa(rom_address_4),
	.datab(rom_address_1),
	.datac(rom_address_0),
	.datad(rom_address_2),
	.cin(gnd),
	.combout(Ram0),
	.cout());
defparam \Ram0~0 .lut_mask = 16'hBFFF;
defparam \Ram0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~3 (
	.dataa(\Ram0~1_combout ),
	.datab(\Ram0~2_combout ),
	.datac(rom_address_4),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Ram01),
	.cout());
defparam \Ram0~3 .lut_mask = 16'h7FF7;
defparam \Ram0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~8 (
	.dataa(Ram0),
	.datab(rom_address_5),
	.datac(\Ram0~6_combout ),
	.datad(\Ram0~7_combout ),
	.cin(gnd),
	.combout(Ram02),
	.cout());
defparam \Ram0~8 .lut_mask = 16'hFFBE;
defparam \Ram0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~9 (
	.dataa(rom_address_0),
	.datab(rom_address_5),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(Ram03),
	.cout());
defparam \Ram0~9 .lut_mask = 16'h6996;
defparam \Ram0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~15 (
	.dataa(\Ram0~10_combout ),
	.datab(rom_address_4),
	.datac(\Ram0~13_combout ),
	.datad(\Ram0~14_combout ),
	.cin(gnd),
	.combout(Ram04),
	.cout());
defparam \Ram0~15 .lut_mask = 16'hFF7D;
defparam \Ram0~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~16 (
	.dataa(rom_address_0),
	.datab(rom_address_4),
	.datac(rom_address_2),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Ram05),
	.cout());
defparam \Ram0~16 .lut_mask = 16'h6996;
defparam \Ram0~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~17 (
	.dataa(rom_address_0),
	.datab(rom_address_4),
	.datac(rom_address_2),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Ram06),
	.cout());
defparam \Ram0~17 .lut_mask = 16'h6996;
defparam \Ram0~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~18 (
	.dataa(rom_address_0),
	.datab(rom_address_4),
	.datac(rom_address_2),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Ram07),
	.cout());
defparam \Ram0~18 .lut_mask = 16'h7FDF;
defparam \Ram0~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~20 (
	.dataa(rom_address_5),
	.datab(\Ram0~19_combout ),
	.datac(rom_address_4),
	.datad(\Ram0~1_combout ),
	.cin(gnd),
	.combout(Ram08),
	.cout());
defparam \Ram0~20 .lut_mask = 16'hFEFF;
defparam \Ram0~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~22 (
	.dataa(rom_address_5),
	.datab(\Ram0~21_combout ),
	.datac(rom_address_4),
	.datad(\Ram0~1_combout ),
	.cin(gnd),
	.combout(Ram09),
	.cout());
defparam \Ram0~22 .lut_mask = 16'hACFF;
defparam \Ram0~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~25 (
	.dataa(\Ram0~24_combout ),
	.datab(rom_address_5),
	.datac(rom_address_4),
	.datad(\Ram0~21_combout ),
	.cin(gnd),
	.combout(Ram010),
	.cout());
defparam \Ram0~25 .lut_mask = 16'hEFFF;
defparam \Ram0~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~1 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~1_combout ),
	.cout());
defparam \Ram0~1 .lut_mask = 16'hFFFE;
defparam \Ram0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~2 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\Ram0~2_combout ),
	.cout());
defparam \Ram0~2 .lut_mask = 16'h7FFF;
defparam \Ram0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~4 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_4),
	.cin(gnd),
	.combout(\Ram0~4_combout ),
	.cout());
defparam \Ram0~4 .lut_mask = 16'hEDDE;
defparam \Ram0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~5 (
	.dataa(rom_address_1),
	.datab(rom_address_4),
	.datac(rom_address_0),
	.datad(rom_address_2),
	.cin(gnd),
	.combout(\Ram0~5_combout ),
	.cout());
defparam \Ram0~5 .lut_mask = 16'hEFFF;
defparam \Ram0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~6 (
	.dataa(rom_address_5),
	.datab(\Ram0~4_combout ),
	.datac(rom_address_3),
	.datad(\Ram0~5_combout ),
	.cin(gnd),
	.combout(\Ram0~6_combout ),
	.cout());
defparam \Ram0~6 .lut_mask = 16'hFFDE;
defparam \Ram0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~7 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_4),
	.cin(gnd),
	.combout(\Ram0~7_combout ),
	.cout());
defparam \Ram0~7 .lut_mask = 16'hF6FF;
defparam \Ram0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~10 (
	.dataa(rom_address_5),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~10_combout ),
	.cout());
defparam \Ram0~10 .lut_mask = 16'hFBFE;
defparam \Ram0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~11 (
	.dataa(rom_address_5),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~11_combout ),
	.cout());
defparam \Ram0~11 .lut_mask = 16'hFFBE;
defparam \Ram0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~12 (
	.dataa(gnd),
	.datab(rom_address_5),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~12_combout ),
	.cout());
defparam \Ram0~12 .lut_mask = 16'hC33C;
defparam \Ram0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~13 (
	.dataa(rom_address_4),
	.datab(\Ram0~11_combout ),
	.datac(rom_address_0),
	.datad(\Ram0~12_combout ),
	.cin(gnd),
	.combout(\Ram0~13_combout ),
	.cout());
defparam \Ram0~13 .lut_mask = 16'hFFDE;
defparam \Ram0~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~14 (
	.dataa(rom_address_5),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~14_combout ),
	.cout());
defparam \Ram0~14 .lut_mask = 16'h6996;
defparam \Ram0~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~19 (
	.dataa(rom_address_2),
	.datab(rom_address_3),
	.datac(gnd),
	.datad(rom_address_4),
	.cin(gnd),
	.combout(\Ram0~19_combout ),
	.cout());
defparam \Ram0~19 .lut_mask = 16'hEEFF;
defparam \Ram0~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~21 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~21_combout ),
	.cout());
defparam \Ram0~21 .lut_mask = 16'hFFFE;
defparam \Ram0~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~23 (
	.dataa(rom_address_0),
	.datab(rom_address_1),
	.datac(rom_address_2),
	.datad(rom_address_3),
	.cin(gnd),
	.combout(\Ram0~23_combout ),
	.cout());
defparam \Ram0~23 .lut_mask = 16'h6996;
defparam \Ram0~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Ram0~24 (
	.dataa(rom_address_4),
	.datab(\Ram0~23_combout ),
	.datac(\Ram0~1_combout ),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(\Ram0~24_combout ),
	.cout());
defparam \Ram0~24 .lut_mask = 16'hFAFC;
defparam \Ram0~24 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_av_config_auto_init_ob_audio (
	rom_address_4,
	rom_address_1,
	rom_address_0,
	rom_address_2,
	rom_address_3,
	rom_address_5,
	Decoder0,
	Decoder01,
	Decoder02,
	Decoder03,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	rom_address_4;
input 	rom_address_1;
input 	rom_address_0;
input 	rom_address_2;
input 	rom_address_3;
input 	rom_address_5;
output 	Decoder0;
output 	Decoder01;
output 	Decoder02;
output 	Decoder03;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \Decoder0~0 (
	.dataa(rom_address_1),
	.datab(rom_address_4),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Decoder0),
	.cout());
defparam \Decoder0~0 .lut_mask = 16'hBFFF;
defparam \Decoder0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~1 (
	.dataa(gnd),
	.datab(rom_address_4),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Decoder01),
	.cout());
defparam \Decoder0~1 .lut_mask = 16'h3FFF;
defparam \Decoder0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~2 (
	.dataa(rom_address_2),
	.datab(rom_address_4),
	.datac(rom_address_3),
	.datad(rom_address_5),
	.cin(gnd),
	.combout(Decoder02),
	.cout());
defparam \Decoder0~2 .lut_mask = 16'hBFFF;
defparam \Decoder0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~3 (
	.dataa(rom_address_0),
	.datab(rom_address_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Decoder03),
	.cout());
defparam \Decoder0~3 .lut_mask = 16'hEEEE;
defparam \Decoder0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(rom_address_1),
	.datab(rom_address_2),
	.datac(rom_address_3),
	.datad(rom_address_4),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hFFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_av_config_serial_bus_controller (
	transfer_data,
	auto_init_complete,
	transfer_complete1,
	shiftreg_data_1,
	shiftreg_data_0,
	shiftreg_data_9,
	shiftreg_data_2,
	shiftreg_data_3,
	shiftreg_data_4,
	shiftreg_data_5,
	data_out_25,
	shiftreg_data_6,
	shiftreg_data_8,
	shiftreg_data_7,
	data_out_1,
	external_read_transfer,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_10,
	data_reg_8,
	data_out_8,
	data_out_7,
	data_out_17,
	data_out_16,
	data_out_15,
	data_out_14,
	data_out_13,
	data_out_12,
	data_out_11,
	serial_clk,
	internal_reset,
	internal_reset1,
	r_sync_rst,
	start_external_transfer,
	shiftreg_mask,
	serial_data,
	serial_data1,
	shiftreg_data_18,
	ack,
	device_for_transfer_1,
	device_for_transfer_0,
	shiftreg_data_10,
	data_reg_0,
	Equal5,
	data_reg_1,
	data_reg_2,
	data_reg_3,
	data_reg_4,
	data_out_24,
	data_reg_5,
	address_for_transfer_0,
	data_reg_7,
	data_reg_6,
	address_for_transfer_7,
	address_for_transfer_6,
	address_for_transfer_5,
	address_for_transfer_4,
	address_for_transfer_3,
	address_for_transfer_2,
	address_for_transfer_1,
	audio_config_wire_SDAT,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	transfer_data;
input 	auto_init_complete;
output 	transfer_complete1;
output 	shiftreg_data_1;
output 	shiftreg_data_0;
output 	shiftreg_data_9;
output 	shiftreg_data_2;
output 	shiftreg_data_3;
output 	shiftreg_data_4;
output 	shiftreg_data_5;
input 	data_out_25;
output 	shiftreg_data_6;
output 	shiftreg_data_8;
output 	shiftreg_data_7;
input 	data_out_1;
input 	external_read_transfer;
input 	data_out_2;
input 	data_out_3;
input 	data_out_4;
input 	data_out_5;
input 	data_out_6;
input 	data_out_10;
input 	data_reg_8;
input 	data_out_8;
input 	data_out_7;
input 	data_out_17;
input 	data_out_16;
input 	data_out_15;
input 	data_out_14;
input 	data_out_13;
input 	data_out_12;
input 	data_out_11;
output 	serial_clk;
input 	internal_reset;
input 	internal_reset1;
input 	r_sync_rst;
input 	start_external_transfer;
output 	shiftreg_mask;
output 	serial_data;
output 	serial_data1;
output 	shiftreg_data_18;
input 	ack;
input 	device_for_transfer_1;
input 	device_for_transfer_0;
output 	shiftreg_data_10;
input 	data_reg_0;
input 	Equal5;
input 	data_reg_1;
input 	data_reg_2;
input 	data_reg_3;
input 	data_reg_4;
input 	data_out_24;
input 	data_reg_5;
input 	address_for_transfer_0;
input 	data_reg_7;
input 	data_reg_6;
input 	address_for_transfer_7;
input 	address_for_transfer_6;
input 	address_for_transfer_5;
input 	address_for_transfer_4;
input 	address_for_transfer_3;
input 	address_for_transfer_2;
input 	address_for_transfer_1;
input 	audio_config_wire_SDAT;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Serial_Config_Clock_Generator|middle_of_high_level~q ;
wire \Serial_Config_Clock_Generator|middle_of_low_level~q ;
wire \Serial_Config_Clock_Generator|new_clk~q ;
wire \Add0~0_combout ;
wire \transfer_complete~0_combout ;
wire \always1~0_combout ;
wire \Selector0~0_combout ;
wire \s_serial_protocol~11_combout ;
wire \s_serial_protocol.STATE_0_IDLE~q ;
wire \s_serial_protocol~12_combout ;
wire \s_serial_protocol.STATE_1_INITIALIZE~q ;
wire \counter~1_combout ;
wire \shiftreg_mask[23]~3_combout ;
wire \shiftreg_mask[23]~4_combout ;
wire \counter[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \Add0~4_combout ;
wire \counter[1]~q ;
wire \Add0~3 ;
wire \Add0~5_combout ;
wire \Add0~9_combout ;
wire \counter[2]~q ;
wire \Add0~6 ;
wire \Add0~7_combout ;
wire \counter~0_combout ;
wire \counter[3]~q ;
wire \always1~1_combout ;
wire \Add0~8 ;
wire \Add0~10_combout ;
wire \Add0~12_combout ;
wire \counter[4]~q ;
wire \Selector1~0_combout ;
wire \shiftreg_data~19_combout ;
wire \shiftreg_data~36_combout ;
wire \shiftreg_data~61_combout ;
wire \shiftreg_data[19]~q ;
wire \shiftreg_data~58_combout ;
wire \shiftreg_data~71_combout ;
wire \shiftreg_data[20]~q ;
wire \shiftreg_data~55_combout ;
wire \shiftreg_data[21]~q ;
wire \shiftreg_data~52_combout ;
wire \shiftreg_data[22]~q ;
wire \shiftreg_data~49_combout ;
wire \shiftreg_data[23]~q ;
wire \shiftreg_data~37_combout ;
wire \shiftreg_data[24]~q ;
wire \shiftreg_data~20_combout ;
wire \shiftreg_data[25]~q ;
wire \shiftreg_data~18_combout ;
wire \shiftreg_data[26]~q ;
wire \shiftreg_mask~31_combout ;
wire \shiftreg_mask[0]~q ;
wire \shiftreg_mask~30_combout ;
wire \shiftreg_mask[1]~q ;
wire \shiftreg_mask~29_combout ;
wire \shiftreg_mask[2]~q ;
wire \shiftreg_mask~28_combout ;
wire \shiftreg_mask[3]~q ;
wire \shiftreg_mask~27_combout ;
wire \shiftreg_mask[4]~q ;
wire \shiftreg_mask~26_combout ;
wire \shiftreg_mask[5]~q ;
wire \shiftreg_mask~25_combout ;
wire \shiftreg_mask[6]~q ;
wire \shiftreg_mask~24_combout ;
wire \shiftreg_mask[7]~q ;
wire \shiftreg_mask~23_combout ;
wire \shiftreg_mask[8]~q ;
wire \shiftreg_mask~22_combout ;
wire \shiftreg_mask[9]~q ;
wire \shiftreg_mask~21_combout ;
wire \shiftreg_mask[10]~q ;
wire \shiftreg_mask~20_combout ;
wire \shiftreg_mask[11]~q ;
wire \shiftreg_mask~19_combout ;
wire \shiftreg_mask[12]~q ;
wire \shiftreg_mask~18_combout ;
wire \shiftreg_mask[13]~q ;
wire \shiftreg_mask~17_combout ;
wire \shiftreg_mask[14]~q ;
wire \shiftreg_mask~16_combout ;
wire \shiftreg_mask[15]~q ;
wire \shiftreg_mask~15_combout ;
wire \shiftreg_mask[16]~q ;
wire \shiftreg_mask~14_combout ;
wire \shiftreg_mask[17]~q ;
wire \shiftreg_mask~13_combout ;
wire \shiftreg_mask[18]~q ;
wire \shiftreg_mask~12_combout ;
wire \shiftreg_mask[19]~q ;
wire \shiftreg_mask~11_combout ;
wire \shiftreg_mask[20]~q ;
wire \shiftreg_mask~10_combout ;
wire \shiftreg_mask[21]~q ;
wire \shiftreg_mask~9_combout ;
wire \shiftreg_mask[22]~q ;
wire \shiftreg_mask~8_combout ;
wire \shiftreg_mask[23]~q ;
wire \shiftreg_mask~7_combout ;
wire \shiftreg_mask[24]~q ;
wire \shiftreg_mask~6_combout ;
wire \shiftreg_mask[25]~q ;
wire \shiftreg_mask~5_combout ;
wire \shiftreg_mask[26]~q ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \s_serial_protocol.STATE_2_RESTART_BIT~q ;
wire \always4~0_combout ;
wire \Selector2~0_combout ;
wire \s_serial_protocol.STATE_3_START_BIT~q ;
wire \Selector3~0_combout ;
wire \s_serial_protocol.STATE_4_TRANSFER~q ;
wire \Selector4~0_combout ;
wire \Selector4~1_combout ;
wire \s_serial_protocol.STATE_5_STOP_BIT~q ;
wire \transfer_complete~1_combout ;
wire \shiftreg_data~21_combout ;
wire \shiftreg_data~22_combout ;
wire \new_data~0_combout ;
wire \new_data~q ;
wire \shiftreg_data~24_combout ;
wire \shiftreg_data~25_combout ;
wire \shiftreg_data[13]~26_combout ;
wire \shiftreg_data~27_combout ;
wire \shiftreg_data~28_combout ;
wire \shiftreg_data~29_combout ;
wire \shiftreg_data~30_combout ;
wire \shiftreg_data~31_combout ;
wire \shiftreg_data~32_combout ;
wire \shiftreg_data~33_combout ;
wire \shiftreg_data~34_combout ;
wire \shiftreg_data~35_combout ;
wire \shiftreg_data~38_combout ;
wire \shiftreg_data~39_combout ;
wire \shiftreg_data~43_combout ;
wire \shiftreg_data~44_combout ;
wire \shiftreg_data~45_combout ;
wire \shiftreg_data~46_combout ;
wire \shiftreg_data[13]~40_combout ;
wire \shiftreg_data~64_combout ;
wire \shiftreg_data~65_combout ;
wire \shiftreg_data~74_combout ;
wire \shiftreg_data[11]~q ;
wire \shiftreg_data~62_combout ;
wire \shiftreg_data~63_combout ;
wire \shiftreg_data~73_combout ;
wire \shiftreg_data[12]~q ;
wire \shiftreg_data~59_combout ;
wire \shiftreg_data~60_combout ;
wire \shiftreg_data~72_combout ;
wire \shiftreg_data[13]~q ;
wire \shiftreg_data~56_combout ;
wire \shiftreg_data~57_combout ;
wire \shiftreg_data~70_combout ;
wire \shiftreg_data[14]~q ;
wire \shiftreg_data~53_combout ;
wire \shiftreg_data~54_combout ;
wire \shiftreg_data~69_combout ;
wire \shiftreg_data[15]~q ;
wire \shiftreg_data~50_combout ;
wire \shiftreg_data~51_combout ;
wire \shiftreg_data~68_combout ;
wire \shiftreg_data[16]~q ;
wire \shiftreg_data~47_combout ;
wire \shiftreg_data~48_combout ;
wire \shiftreg_data~67_combout ;
wire \shiftreg_data[17]~q ;
wire \shiftreg_data~23_combout ;
wire \shiftreg_data~41_combout ;
wire \shiftreg_data~42_combout ;
wire \shiftreg_data~66_combout ;


final_project_soc_altera_up_slow_clock_generator Serial_Config_Clock_Generator(
	.middle_of_high_level1(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.middle_of_low_level1(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.new_clk1(\Serial_Config_Clock_Generator|new_clk~q ),
	.internal_reset(internal_reset),
	.internal_reset1(internal_reset1),
	.r_sync_rst(r_sync_rst),
	.shiftreg_mask(shiftreg_mask),
	.clk(clk_clk));

dffeas transfer_complete(
	.clk(clk_clk),
	.d(\transfer_complete~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(transfer_complete1),
	.prn(vcc));
defparam transfer_complete.is_wysiwyg = "true";
defparam transfer_complete.power_up = "low";

dffeas \shiftreg_data[1] (
	.clk(clk_clk),
	.d(\shiftreg_data~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_1),
	.prn(vcc));
defparam \shiftreg_data[1] .is_wysiwyg = "true";
defparam \shiftreg_data[1] .power_up = "low";

dffeas \shiftreg_data[0] (
	.clk(clk_clk),
	.d(\shiftreg_data~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_0),
	.prn(vcc));
defparam \shiftreg_data[0] .is_wysiwyg = "true";
defparam \shiftreg_data[0] .power_up = "low";

dffeas \shiftreg_data[9] (
	.clk(clk_clk),
	.d(\shiftreg_data~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_9),
	.prn(vcc));
defparam \shiftreg_data[9] .is_wysiwyg = "true";
defparam \shiftreg_data[9] .power_up = "low";

dffeas \shiftreg_data[2] (
	.clk(clk_clk),
	.d(\shiftreg_data~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_2),
	.prn(vcc));
defparam \shiftreg_data[2] .is_wysiwyg = "true";
defparam \shiftreg_data[2] .power_up = "low";

dffeas \shiftreg_data[3] (
	.clk(clk_clk),
	.d(\shiftreg_data~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_3),
	.prn(vcc));
defparam \shiftreg_data[3] .is_wysiwyg = "true";
defparam \shiftreg_data[3] .power_up = "low";

dffeas \shiftreg_data[4] (
	.clk(clk_clk),
	.d(\shiftreg_data~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_4),
	.prn(vcc));
defparam \shiftreg_data[4] .is_wysiwyg = "true";
defparam \shiftreg_data[4] .power_up = "low";

dffeas \shiftreg_data[5] (
	.clk(clk_clk),
	.d(\shiftreg_data~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_5),
	.prn(vcc));
defparam \shiftreg_data[5] .is_wysiwyg = "true";
defparam \shiftreg_data[5] .power_up = "low";

dffeas \shiftreg_data[6] (
	.clk(clk_clk),
	.d(\shiftreg_data~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_6),
	.prn(vcc));
defparam \shiftreg_data[6] .is_wysiwyg = "true";
defparam \shiftreg_data[6] .power_up = "low";

dffeas \shiftreg_data[8] (
	.clk(clk_clk),
	.d(\shiftreg_data~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_8),
	.prn(vcc));
defparam \shiftreg_data[8] .is_wysiwyg = "true";
defparam \shiftreg_data[8] .power_up = "low";

dffeas \shiftreg_data[7] (
	.clk(clk_clk),
	.d(\shiftreg_data~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_7),
	.prn(vcc));
defparam \shiftreg_data[7] .is_wysiwyg = "true";
defparam \shiftreg_data[7] .power_up = "low";

cycloneive_lcell_comb \serial_clk~0 (
	.dataa(\Serial_Config_Clock_Generator|new_clk~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\s_serial_protocol.STATE_0_IDLE~q ),
	.cin(gnd),
	.combout(serial_clk),
	.cout());
defparam \serial_clk~0 .lut_mask = 16'hAAFF;
defparam \serial_clk~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_mask~2 (
	.dataa(gnd),
	.datab(internal_reset),
	.datac(internal_reset1),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(shiftreg_mask),
	.cout());
defparam \shiftreg_mask~2 .lut_mask = 16'hFFFC;
defparam \shiftreg_mask~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \serial_data~1 (
	.dataa(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datab(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.datac(\shiftreg_data[26]~q ),
	.datad(\s_serial_protocol.STATE_0_IDLE~q ),
	.cin(gnd),
	.combout(serial_data),
	.cout());
defparam \serial_data~1 .lut_mask = 16'hFEFF;
defparam \serial_data~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \serial_data~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.datad(\shiftreg_mask[26]~q ),
	.cin(gnd),
	.combout(serial_data1),
	.cout());
defparam \serial_data~2 .lut_mask = 16'h0FFF;
defparam \serial_data~2 .sum_lutc_input = "datac";

dffeas \shiftreg_data[18] (
	.clk(clk_clk),
	.d(\shiftreg_data~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_18),
	.prn(vcc));
defparam \shiftreg_data[18] .is_wysiwyg = "true";
defparam \shiftreg_data[18] .power_up = "low";

dffeas \shiftreg_data[10] (
	.clk(clk_clk),
	.d(\shiftreg_data~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(shiftreg_data_10),
	.prn(vcc));
defparam \shiftreg_data[10] .is_wysiwyg = "true";
defparam \shiftreg_data[10] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \transfer_complete~0 (
	.dataa(start_external_transfer),
	.datab(transfer_data),
	.datac(gnd),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\transfer_complete~0_combout ),
	.cout());
defparam \transfer_complete~0 .lut_mask = 16'hAACC;
defparam \transfer_complete~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\transfer_complete~0_combout ),
	.datac(gnd),
	.datad(transfer_complete1),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hEEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_5_STOP_BIT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEEEE;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \s_serial_protocol~11 (
	.dataa(\Selector0~0_combout ),
	.datab(\s_serial_protocol.STATE_0_IDLE~q ),
	.datac(\always1~0_combout ),
	.datad(shiftreg_mask),
	.cin(gnd),
	.combout(\s_serial_protocol~11_combout ),
	.cout());
defparam \s_serial_protocol~11 .lut_mask = 16'hFDFF;
defparam \s_serial_protocol~11 .sum_lutc_input = "datac";

dffeas \s_serial_protocol.STATE_0_IDLE (
	.clk(clk_clk),
	.d(\s_serial_protocol~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_protocol.STATE_0_IDLE~q ),
	.prn(vcc));
defparam \s_serial_protocol.STATE_0_IDLE .is_wysiwyg = "true";
defparam \s_serial_protocol.STATE_0_IDLE .power_up = "low";

cycloneive_lcell_comb \s_serial_protocol~12 (
	.dataa(shiftreg_mask),
	.datab(\always1~0_combout ),
	.datac(gnd),
	.datad(\s_serial_protocol.STATE_0_IDLE~q ),
	.cin(gnd),
	.combout(\s_serial_protocol~12_combout ),
	.cout());
defparam \s_serial_protocol~12 .lut_mask = 16'hDDFF;
defparam \s_serial_protocol~12 .sum_lutc_input = "datac";

dffeas \s_serial_protocol.STATE_1_INITIALIZE (
	.clk(clk_clk),
	.d(\s_serial_protocol~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.prn(vcc));
defparam \s_serial_protocol.STATE_1_INITIALIZE .is_wysiwyg = "true";
defparam \s_serial_protocol.STATE_1_INITIALIZE .power_up = "low";

cycloneive_lcell_comb \counter~1 (
	.dataa(shiftreg_mask),
	.datab(\Add0~0_combout ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\counter~1_combout ),
	.cout());
defparam \counter~1 .lut_mask = 16'hFDFF;
defparam \counter~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_mask[23]~3 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(r_sync_rst),
	.datac(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.datad(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.cin(gnd),
	.combout(\shiftreg_mask[23]~3_combout ),
	.cout());
defparam \shiftreg_mask[23]~3 .lut_mask = 16'hFFFE;
defparam \shiftreg_mask[23]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_mask[23]~4 (
	.dataa(\always4~0_combout ),
	.datab(internal_reset),
	.datac(internal_reset1),
	.datad(\shiftreg_mask[23]~3_combout ),
	.cin(gnd),
	.combout(\shiftreg_mask[23]~4_combout ),
	.cout());
defparam \shiftreg_mask[23]~4 .lut_mask = 16'hFFFE;
defparam \shiftreg_mask[23]~4 .sum_lutc_input = "datac";

dffeas \counter[0] (
	.clk(clk_clk),
	.d(\counter~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\counter[0]~q ),
	.prn(vcc));
defparam \counter[0] .is_wysiwyg = "true";
defparam \counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(shiftreg_mask),
	.datab(\Add0~2_combout ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\Add0~4_combout ),
	.cout());
defparam \Add0~4 .lut_mask = 16'hDFFF;
defparam \Add0~4 .sum_lutc_input = "datac";

dffeas \counter[1] (
	.clk(clk_clk),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\counter[1]~q ),
	.prn(vcc));
defparam \counter[1] .is_wysiwyg = "true";
defparam \counter[1] .power_up = "low";

cycloneive_lcell_comb \Add0~5 (
	.dataa(\counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~5_combout ),
	.cout(\Add0~6 ));
defparam \Add0~5 .lut_mask = 16'h5AAF;
defparam \Add0~5 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~9 (
	.dataa(shiftreg_mask),
	.datab(\Add0~5_combout ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\Add0~9_combout ),
	.cout());
defparam \Add0~9 .lut_mask = 16'hDFFF;
defparam \Add0~9 .sum_lutc_input = "datac";

dffeas \counter[2] (
	.clk(clk_clk),
	.d(\Add0~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\counter[2]~q ),
	.prn(vcc));
defparam \counter[2] .is_wysiwyg = "true";
defparam \counter[2] .power_up = "low";

cycloneive_lcell_comb \Add0~7 (
	.dataa(\counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~6 ),
	.combout(\Add0~7_combout ),
	.cout(\Add0~8 ));
defparam \Add0~7 .lut_mask = 16'h5A5F;
defparam \Add0~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \counter~0 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\Add0~7_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\counter~0_combout ),
	.cout());
defparam \counter~0 .lut_mask = 16'hFDFF;
defparam \counter~0 .sum_lutc_input = "datac";

dffeas \counter[3] (
	.clk(clk_clk),
	.d(\counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\counter[3]~q ),
	.prn(vcc));
defparam \counter[3] .is_wysiwyg = "true";
defparam \counter[3] .power_up = "low";

cycloneive_lcell_comb \always1~1 (
	.dataa(\counter[1]~q ),
	.datab(\counter[3]~q ),
	.datac(\counter[0]~q ),
	.datad(\counter[2]~q ),
	.cin(gnd),
	.combout(\always1~1_combout ),
	.cout());
defparam \always1~1 .lut_mask = 16'hEFFF;
defparam \always1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~10 (
	.dataa(\counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~8 ),
	.combout(\Add0~10_combout ),
	.cout());
defparam \Add0~10 .lut_mask = 16'h5A5A;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~12 (
	.dataa(shiftreg_mask),
	.datab(\Add0~10_combout ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'hDFFF;
defparam \Add0~12 .sum_lutc_input = "datac";

dffeas \counter[4] (
	.clk(clk_clk),
	.d(\Add0~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\counter[4]~q ),
	.prn(vcc));
defparam \counter[4] .is_wysiwyg = "true";
defparam \counter[4] .power_up = "low";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.datab(\always1~1_combout ),
	.datac(\counter[4]~q ),
	.datad(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hBFFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~19 (
	.dataa(data_out_25),
	.datab(auto_init_complete),
	.datac(device_for_transfer_1),
	.datad(device_for_transfer_0),
	.cin(gnd),
	.combout(\shiftreg_data~19_combout ),
	.cout());
defparam \shiftreg_data~19 .lut_mask = 16'hFFB8;
defparam \shiftreg_data~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~36 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_out_24),
	.datac(auto_init_complete),
	.datad(Equal5),
	.cin(gnd),
	.combout(\shiftreg_data~36_combout ),
	.cout());
defparam \shiftreg_data~36 .lut_mask = 16'hACFF;
defparam \shiftreg_data~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~61 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(shiftreg_data_18),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~61_combout ),
	.cout());
defparam \shiftreg_data~61 .lut_mask = 16'hFDFF;
defparam \shiftreg_data~61 .sum_lutc_input = "datac";

dffeas \shiftreg_data[19] (
	.clk(clk_clk),
	.d(\shiftreg_data~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[19]~q ),
	.prn(vcc));
defparam \shiftreg_data[19] .is_wysiwyg = "true";
defparam \shiftreg_data[19] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~58 (
	.dataa(device_for_transfer_1),
	.datab(\shiftreg_data[19]~q ),
	.datac(\always4~0_combout ),
	.datad(device_for_transfer_0),
	.cin(gnd),
	.combout(\shiftreg_data~58_combout ),
	.cout());
defparam \shiftreg_data~58 .lut_mask = 16'hACFF;
defparam \shiftreg_data~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~71 (
	.dataa(auto_init_complete),
	.datab(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datac(device_for_transfer_1),
	.datad(\shiftreg_data~58_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~71_combout ),
	.cout());
defparam \shiftreg_data~71 .lut_mask = 16'hFFB8;
defparam \shiftreg_data~71 .sum_lutc_input = "datac";

dffeas \shiftreg_data[20] (
	.clk(clk_clk),
	.d(\shiftreg_data~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[20]~q ),
	.prn(vcc));
defparam \shiftreg_data[20] .is_wysiwyg = "true";
defparam \shiftreg_data[20] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~55 (
	.dataa(\shiftreg_data~36_combout ),
	.datab(\shiftreg_data[20]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~55_combout ),
	.cout());
defparam \shiftreg_data~55 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~55 .sum_lutc_input = "datac";

dffeas \shiftreg_data[21] (
	.clk(clk_clk),
	.d(\shiftreg_data~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[21]~q ),
	.prn(vcc));
defparam \shiftreg_data[21] .is_wysiwyg = "true";
defparam \shiftreg_data[21] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~52 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_data[21]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~52_combout ),
	.cout());
defparam \shiftreg_data~52 .lut_mask = 16'hDFFF;
defparam \shiftreg_data~52 .sum_lutc_input = "datac";

dffeas \shiftreg_data[22] (
	.clk(clk_clk),
	.d(\shiftreg_data~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[22]~q ),
	.prn(vcc));
defparam \shiftreg_data[22] .is_wysiwyg = "true";
defparam \shiftreg_data[22] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~49 (
	.dataa(\shiftreg_data~36_combout ),
	.datab(\shiftreg_data[22]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~49_combout ),
	.cout());
defparam \shiftreg_data~49 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~49 .sum_lutc_input = "datac";

dffeas \shiftreg_data[23] (
	.clk(clk_clk),
	.d(\shiftreg_data~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[23]~q ),
	.prn(vcc));
defparam \shiftreg_data[23] .is_wysiwyg = "true";
defparam \shiftreg_data[23] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~37 (
	.dataa(\shiftreg_data~36_combout ),
	.datab(\shiftreg_data[23]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~37_combout ),
	.cout());
defparam \shiftreg_data~37 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~37 .sum_lutc_input = "datac";

dffeas \shiftreg_data[24] (
	.clk(clk_clk),
	.d(\shiftreg_data~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[24]~q ),
	.prn(vcc));
defparam \shiftreg_data[24] .is_wysiwyg = "true";
defparam \shiftreg_data[24] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~20 (
	.dataa(\shiftreg_data~19_combout ),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_data[24]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~20_combout ),
	.cout());
defparam \shiftreg_data~20 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~20 .sum_lutc_input = "datac";

dffeas \shiftreg_data[25] (
	.clk(clk_clk),
	.d(\shiftreg_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[25]~q ),
	.prn(vcc));
defparam \shiftreg_data[25] .is_wysiwyg = "true";
defparam \shiftreg_data[25] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~18 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_data[25]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~18_combout ),
	.cout());
defparam \shiftreg_data~18 .lut_mask = 16'hDFFF;
defparam \shiftreg_data~18 .sum_lutc_input = "datac";

dffeas \shiftreg_data[26] (
	.clk(clk_clk),
	.d(\shiftreg_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[26]~q ),
	.prn(vcc));
defparam \shiftreg_data[26] .is_wysiwyg = "true";
defparam \shiftreg_data[26] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~31 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~31_combout ),
	.cout());
defparam \shiftreg_mask~31 .lut_mask = 16'hFFEF;
defparam \shiftreg_mask~31 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[0] (
	.clk(clk_clk),
	.d(\shiftreg_mask~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[0]~q ),
	.prn(vcc));
defparam \shiftreg_mask[0] .is_wysiwyg = "true";
defparam \shiftreg_mask[0] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~30 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[0]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~30_combout ),
	.cout());
defparam \shiftreg_mask~30 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~30 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[1] (
	.clk(clk_clk),
	.d(\shiftreg_mask~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[1]~q ),
	.prn(vcc));
defparam \shiftreg_mask[1] .is_wysiwyg = "true";
defparam \shiftreg_mask[1] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~29 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[1]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~29_combout ),
	.cout());
defparam \shiftreg_mask~29 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~29 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[2] (
	.clk(clk_clk),
	.d(\shiftreg_mask~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[2]~q ),
	.prn(vcc));
defparam \shiftreg_mask[2] .is_wysiwyg = "true";
defparam \shiftreg_mask[2] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~28 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[2]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~28_combout ),
	.cout());
defparam \shiftreg_mask~28 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~28 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[3] (
	.clk(clk_clk),
	.d(\shiftreg_mask~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[3]~q ),
	.prn(vcc));
defparam \shiftreg_mask[3] .is_wysiwyg = "true";
defparam \shiftreg_mask[3] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~27 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[3]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~27_combout ),
	.cout());
defparam \shiftreg_mask~27 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~27 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[4] (
	.clk(clk_clk),
	.d(\shiftreg_mask~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[4]~q ),
	.prn(vcc));
defparam \shiftreg_mask[4] .is_wysiwyg = "true";
defparam \shiftreg_mask[4] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~26 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[4]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~26_combout ),
	.cout());
defparam \shiftreg_mask~26 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~26 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[5] (
	.clk(clk_clk),
	.d(\shiftreg_mask~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[5]~q ),
	.prn(vcc));
defparam \shiftreg_mask[5] .is_wysiwyg = "true";
defparam \shiftreg_mask[5] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~25 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[5]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~25_combout ),
	.cout());
defparam \shiftreg_mask~25 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~25 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[6] (
	.clk(clk_clk),
	.d(\shiftreg_mask~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[6]~q ),
	.prn(vcc));
defparam \shiftreg_mask[6] .is_wysiwyg = "true";
defparam \shiftreg_mask[6] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~24 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[6]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~24_combout ),
	.cout());
defparam \shiftreg_mask~24 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~24 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[7] (
	.clk(clk_clk),
	.d(\shiftreg_mask~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[7]~q ),
	.prn(vcc));
defparam \shiftreg_mask[7] .is_wysiwyg = "true";
defparam \shiftreg_mask[7] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~23 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[7]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~23_combout ),
	.cout());
defparam \shiftreg_mask~23 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~23 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[8] (
	.clk(clk_clk),
	.d(\shiftreg_mask~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[8]~q ),
	.prn(vcc));
defparam \shiftreg_mask[8] .is_wysiwyg = "true";
defparam \shiftreg_mask[8] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~22 (
	.dataa(shiftreg_mask),
	.datab(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datac(\shiftreg_mask[8]~q ),
	.datad(\always4~0_combout ),
	.cin(gnd),
	.combout(\shiftreg_mask~22_combout ),
	.cout());
defparam \shiftreg_mask~22 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~22 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[9] (
	.clk(clk_clk),
	.d(\shiftreg_mask~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[9]~q ),
	.prn(vcc));
defparam \shiftreg_mask[9] .is_wysiwyg = "true";
defparam \shiftreg_mask[9] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~21 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[9]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~21_combout ),
	.cout());
defparam \shiftreg_mask~21 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~21 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[10] (
	.clk(clk_clk),
	.d(\shiftreg_mask~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[10]~q ),
	.prn(vcc));
defparam \shiftreg_mask[10] .is_wysiwyg = "true";
defparam \shiftreg_mask[10] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~20 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[10]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~20_combout ),
	.cout());
defparam \shiftreg_mask~20 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~20 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[11] (
	.clk(clk_clk),
	.d(\shiftreg_mask~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[11]~q ),
	.prn(vcc));
defparam \shiftreg_mask[11] .is_wysiwyg = "true";
defparam \shiftreg_mask[11] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~19 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[11]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~19_combout ),
	.cout());
defparam \shiftreg_mask~19 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~19 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[12] (
	.clk(clk_clk),
	.d(\shiftreg_mask~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[12]~q ),
	.prn(vcc));
defparam \shiftreg_mask[12] .is_wysiwyg = "true";
defparam \shiftreg_mask[12] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~18 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[12]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~18_combout ),
	.cout());
defparam \shiftreg_mask~18 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~18 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[13] (
	.clk(clk_clk),
	.d(\shiftreg_mask~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[13]~q ),
	.prn(vcc));
defparam \shiftreg_mask[13] .is_wysiwyg = "true";
defparam \shiftreg_mask[13] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~17 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[13]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~17_combout ),
	.cout());
defparam \shiftreg_mask~17 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~17 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[14] (
	.clk(clk_clk),
	.d(\shiftreg_mask~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[14]~q ),
	.prn(vcc));
defparam \shiftreg_mask[14] .is_wysiwyg = "true";
defparam \shiftreg_mask[14] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~16 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[14]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~16_combout ),
	.cout());
defparam \shiftreg_mask~16 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~16 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[15] (
	.clk(clk_clk),
	.d(\shiftreg_mask~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[15]~q ),
	.prn(vcc));
defparam \shiftreg_mask[15] .is_wysiwyg = "true";
defparam \shiftreg_mask[15] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~15 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[15]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~15_combout ),
	.cout());
defparam \shiftreg_mask~15 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~15 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[16] (
	.clk(clk_clk),
	.d(\shiftreg_mask~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[16]~q ),
	.prn(vcc));
defparam \shiftreg_mask[16] .is_wysiwyg = "true";
defparam \shiftreg_mask[16] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~14 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\shiftreg_mask[16]~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~14_combout ),
	.cout());
defparam \shiftreg_mask~14 .lut_mask = 16'hFDFF;
defparam \shiftreg_mask~14 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[17] (
	.clk(clk_clk),
	.d(\shiftreg_mask~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[17]~q ),
	.prn(vcc));
defparam \shiftreg_mask[17] .is_wysiwyg = "true";
defparam \shiftreg_mask[17] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~13 (
	.dataa(shiftreg_mask),
	.datab(\always4~0_combout ),
	.datac(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datad(\shiftreg_mask[17]~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~13_combout ),
	.cout());
defparam \shiftreg_mask~13 .lut_mask = 16'hFFFD;
defparam \shiftreg_mask~13 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[18] (
	.clk(clk_clk),
	.d(\shiftreg_mask~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[18]~q ),
	.prn(vcc));
defparam \shiftreg_mask[18] .is_wysiwyg = "true";
defparam \shiftreg_mask[18] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~12 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[18]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~12_combout ),
	.cout());
defparam \shiftreg_mask~12 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~12 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[19] (
	.clk(clk_clk),
	.d(\shiftreg_mask~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[19]~q ),
	.prn(vcc));
defparam \shiftreg_mask[19] .is_wysiwyg = "true";
defparam \shiftreg_mask[19] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~11 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[19]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~11_combout ),
	.cout());
defparam \shiftreg_mask~11 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~11 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[20] (
	.clk(clk_clk),
	.d(\shiftreg_mask~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[20]~q ),
	.prn(vcc));
defparam \shiftreg_mask[20] .is_wysiwyg = "true";
defparam \shiftreg_mask[20] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~10 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[20]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~10_combout ),
	.cout());
defparam \shiftreg_mask~10 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~10 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[21] (
	.clk(clk_clk),
	.d(\shiftreg_mask~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[21]~q ),
	.prn(vcc));
defparam \shiftreg_mask[21] .is_wysiwyg = "true";
defparam \shiftreg_mask[21] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~9 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[21]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~9_combout ),
	.cout());
defparam \shiftreg_mask~9 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~9 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[22] (
	.clk(clk_clk),
	.d(\shiftreg_mask~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[22]~q ),
	.prn(vcc));
defparam \shiftreg_mask[22] .is_wysiwyg = "true";
defparam \shiftreg_mask[22] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~8 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[22]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~8_combout ),
	.cout());
defparam \shiftreg_mask~8 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~8 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[23] (
	.clk(clk_clk),
	.d(\shiftreg_mask~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[23]~q ),
	.prn(vcc));
defparam \shiftreg_mask[23] .is_wysiwyg = "true";
defparam \shiftreg_mask[23] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~7 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[23]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~7_combout ),
	.cout());
defparam \shiftreg_mask~7 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~7 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[24] (
	.clk(clk_clk),
	.d(\shiftreg_mask~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[24]~q ),
	.prn(vcc));
defparam \shiftreg_mask[24] .is_wysiwyg = "true";
defparam \shiftreg_mask[24] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~6 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[24]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~6_combout ),
	.cout());
defparam \shiftreg_mask~6 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~6 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[25] (
	.clk(clk_clk),
	.d(\shiftreg_mask~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[25]~q ),
	.prn(vcc));
defparam \shiftreg_mask[25] .is_wysiwyg = "true";
defparam \shiftreg_mask[25] .power_up = "low";

cycloneive_lcell_comb \shiftreg_mask~5 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_mask[25]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_mask~5_combout ),
	.cout());
defparam \shiftreg_mask~5 .lut_mask = 16'hDFFF;
defparam \shiftreg_mask~5 .sum_lutc_input = "datac";

dffeas \shiftreg_mask[26] (
	.clk(clk_clk),
	.d(\shiftreg_mask~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_mask[26]~q ),
	.prn(vcc));
defparam \shiftreg_mask[26] .is_wysiwyg = "true";
defparam \shiftreg_mask[26] .power_up = "low";

cycloneive_lcell_comb \Selector1~1 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.datab(\shiftreg_data[26]~q ),
	.datac(\shiftreg_mask[26]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hFEFE;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datad(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFEFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \s_serial_protocol.STATE_2_RESTART_BIT (
	.clk(clk_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.prn(vcc));
defparam \s_serial_protocol.STATE_2_RESTART_BIT .is_wysiwyg = "true";
defparam \s_serial_protocol.STATE_2_RESTART_BIT .power_up = "low";

cycloneive_lcell_comb \always4~0 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hEEEE;
defparam \always4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\always4~0_combout ),
	.datab(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datac(\s_serial_protocol.STATE_3_START_BIT~q ),
	.datad(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \s_serial_protocol.STATE_3_START_BIT (
	.clk(clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_protocol.STATE_3_START_BIT~q ),
	.prn(vcc));
defparam \s_serial_protocol.STATE_3_START_BIT .is_wysiwyg = "true";
defparam \s_serial_protocol.STATE_3_START_BIT .power_up = "low";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.datab(\s_serial_protocol.STATE_3_START_BIT~q ),
	.datac(\Selector1~0_combout ),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFEFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \s_serial_protocol.STATE_4_TRANSFER (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.prn(vcc));
defparam \s_serial_protocol.STATE_4_TRANSFER .is_wysiwyg = "true";
defparam \s_serial_protocol.STATE_4_TRANSFER .power_up = "low";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.datab(\always1~1_combout ),
	.datac(\counter[4]~q ),
	.datad(\Serial_Config_Clock_Generator|middle_of_low_level~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFFFE;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(\Selector4~0_combout ),
	.datab(\s_serial_protocol.STATE_5_STOP_BIT~q ),
	.datac(gnd),
	.datad(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hEEFF;
defparam \Selector4~1 .sum_lutc_input = "datac";

dffeas \s_serial_protocol.STATE_5_STOP_BIT (
	.clk(clk_clk),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\s_serial_protocol.STATE_5_STOP_BIT~q ),
	.prn(vcc));
defparam \s_serial_protocol.STATE_5_STOP_BIT .is_wysiwyg = "true";
defparam \s_serial_protocol.STATE_5_STOP_BIT .power_up = "low";

cycloneive_lcell_comb \transfer_complete~1 (
	.dataa(\s_serial_protocol.STATE_5_STOP_BIT~q ),
	.datab(transfer_complete1),
	.datac(\transfer_complete~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\transfer_complete~1_combout ),
	.cout());
defparam \transfer_complete~1 .lut_mask = 16'hFEFE;
defparam \transfer_complete~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~21 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_0),
	.datac(data_out_1),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~21_combout ),
	.cout());
defparam \shiftreg_data~21 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~22 (
	.dataa(\shiftreg_data~21_combout ),
	.datab(shiftreg_data_0),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~22_combout ),
	.cout());
defparam \shiftreg_data~22 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \new_data~0 (
	.dataa(audio_config_wire_SDAT),
	.datab(\new_data~q ),
	.datac(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datad(\s_serial_protocol.STATE_4_TRANSFER~q ),
	.cin(gnd),
	.combout(\new_data~0_combout ),
	.cout());
defparam \new_data~0 .lut_mask = 16'hEFFE;
defparam \new_data~0 .sum_lutc_input = "datac";

dffeas new_data(
	.clk(clk_clk),
	.d(\new_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\new_data~q ),
	.prn(vcc));
defparam new_data.is_wysiwyg = "true";
defparam new_data.power_up = "low";

cycloneive_lcell_comb \shiftreg_data~24 (
	.dataa(shiftreg_mask),
	.datab(ack),
	.datac(\new_data~q ),
	.datad(\always4~0_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~24_combout ),
	.cout());
defparam \shiftreg_data~24 .lut_mask = 16'hDDF5;
defparam \shiftreg_data~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~25 (
	.dataa(shiftreg_data_8),
	.datab(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datac(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~25_combout ),
	.cout());
defparam \shiftreg_data~25 .lut_mask = 16'hBFFF;
defparam \shiftreg_data~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data[13]~26 (
	.dataa(auto_init_complete),
	.datab(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\shiftreg_data[13]~26_combout ),
	.cout());
defparam \shiftreg_data[13]~26 .lut_mask = 16'hEEEE;
defparam \shiftreg_data[13]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~27 (
	.dataa(\shiftreg_data~25_combout ),
	.datab(Equal5),
	.datac(external_read_transfer),
	.datad(\shiftreg_data[13]~26_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~27_combout ),
	.cout());
defparam \shiftreg_data~27 .lut_mask = 16'hFFFE;
defparam \shiftreg_data~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~28 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_1),
	.datac(data_out_2),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~28_combout ),
	.cout());
defparam \shiftreg_data~28 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~29 (
	.dataa(\shiftreg_data~28_combout ),
	.datab(shiftreg_data_1),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~29_combout ),
	.cout());
defparam \shiftreg_data~29 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~30 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_2),
	.datac(data_out_3),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~30_combout ),
	.cout());
defparam \shiftreg_data~30 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~31 (
	.dataa(\shiftreg_data~30_combout ),
	.datab(shiftreg_data_2),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~31_combout ),
	.cout());
defparam \shiftreg_data~31 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~32 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_3),
	.datac(data_out_4),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~32_combout ),
	.cout());
defparam \shiftreg_data~32 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~33 (
	.dataa(\shiftreg_data~32_combout ),
	.datab(shiftreg_data_3),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~33_combout ),
	.cout());
defparam \shiftreg_data~33 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~34 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_4),
	.datac(data_out_5),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~34_combout ),
	.cout());
defparam \shiftreg_data~34 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~35 (
	.dataa(\shiftreg_data~34_combout ),
	.datab(shiftreg_data_4),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~35_combout ),
	.cout());
defparam \shiftreg_data~35 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~38 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_5),
	.datac(data_out_6),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~38_combout ),
	.cout());
defparam \shiftreg_data~38 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~39 (
	.dataa(\shiftreg_data~38_combout ),
	.datab(shiftreg_data_5),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~39_combout ),
	.cout());
defparam \shiftreg_data~39 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~43 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_7),
	.datac(data_out_8),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~43_combout ),
	.cout());
defparam \shiftreg_data~43 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~44 (
	.dataa(\shiftreg_data~43_combout ),
	.datab(shiftreg_data_7),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~44_combout ),
	.cout());
defparam \shiftreg_data~44 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~45 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(data_reg_6),
	.datac(data_out_7),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data~45_combout ),
	.cout());
defparam \shiftreg_data~45 .lut_mask = 16'hFAFC;
defparam \shiftreg_data~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~46 (
	.dataa(\shiftreg_data~45_combout ),
	.datab(shiftreg_data_6),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~46_combout ),
	.cout());
defparam \shiftreg_data~46 .lut_mask = 16'hEFFF;
defparam \shiftreg_data~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data[13]~40 (
	.dataa(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.datab(device_for_transfer_1),
	.datac(device_for_transfer_0),
	.datad(auto_init_complete),
	.cin(gnd),
	.combout(\shiftreg_data[13]~40_combout ),
	.cout());
defparam \shiftreg_data[13]~40 .lut_mask = 16'hBFFF;
defparam \shiftreg_data[13]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~64 (
	.dataa(\shiftreg_data[13]~26_combout ),
	.datab(data_out_11),
	.datac(\shiftreg_data[13]~40_combout ),
	.datad(shiftreg_data_10),
	.cin(gnd),
	.combout(\shiftreg_data~64_combout ),
	.cout());
defparam \shiftreg_data~64 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~65 (
	.dataa(address_for_transfer_1),
	.datab(\shiftreg_data[13]~26_combout ),
	.datac(\shiftreg_data~64_combout ),
	.datad(address_for_transfer_0),
	.cin(gnd),
	.combout(\shiftreg_data~65_combout ),
	.cout());
defparam \shiftreg_data~65 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~74 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~65_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~74_combout ),
	.cout());
defparam \shiftreg_data~74 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~74 .sum_lutc_input = "datac";

dffeas \shiftreg_data[11] (
	.clk(clk_clk),
	.d(\shiftreg_data~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[11]~q ),
	.prn(vcc));
defparam \shiftreg_data[11] .is_wysiwyg = "true";
defparam \shiftreg_data[11] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~62 (
	.dataa(\shiftreg_data[13]~40_combout ),
	.datab(address_for_transfer_2),
	.datac(\shiftreg_data[13]~26_combout ),
	.datad(\shiftreg_data[11]~q ),
	.cin(gnd),
	.combout(\shiftreg_data~62_combout ),
	.cout());
defparam \shiftreg_data~62 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~63 (
	.dataa(data_out_12),
	.datab(\shiftreg_data[13]~40_combout ),
	.datac(\shiftreg_data~62_combout ),
	.datad(address_for_transfer_1),
	.cin(gnd),
	.combout(\shiftreg_data~63_combout ),
	.cout());
defparam \shiftreg_data~63 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~73 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~63_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~73_combout ),
	.cout());
defparam \shiftreg_data~73 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~73 .sum_lutc_input = "datac";

dffeas \shiftreg_data[12] (
	.clk(clk_clk),
	.d(\shiftreg_data~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[12]~q ),
	.prn(vcc));
defparam \shiftreg_data[12] .is_wysiwyg = "true";
defparam \shiftreg_data[12] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~59 (
	.dataa(\shiftreg_data[13]~26_combout ),
	.datab(data_out_13),
	.datac(\shiftreg_data[13]~40_combout ),
	.datad(\shiftreg_data[12]~q ),
	.cin(gnd),
	.combout(\shiftreg_data~59_combout ),
	.cout());
defparam \shiftreg_data~59 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~60 (
	.dataa(address_for_transfer_3),
	.datab(\shiftreg_data[13]~26_combout ),
	.datac(\shiftreg_data~59_combout ),
	.datad(address_for_transfer_2),
	.cin(gnd),
	.combout(\shiftreg_data~60_combout ),
	.cout());
defparam \shiftreg_data~60 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~72 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~60_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~72_combout ),
	.cout());
defparam \shiftreg_data~72 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~72 .sum_lutc_input = "datac";

dffeas \shiftreg_data[13] (
	.clk(clk_clk),
	.d(\shiftreg_data~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[13]~q ),
	.prn(vcc));
defparam \shiftreg_data[13] .is_wysiwyg = "true";
defparam \shiftreg_data[13] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~56 (
	.dataa(\shiftreg_data[13]~40_combout ),
	.datab(address_for_transfer_4),
	.datac(\shiftreg_data[13]~26_combout ),
	.datad(\shiftreg_data[13]~q ),
	.cin(gnd),
	.combout(\shiftreg_data~56_combout ),
	.cout());
defparam \shiftreg_data~56 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~57 (
	.dataa(data_out_14),
	.datab(\shiftreg_data[13]~40_combout ),
	.datac(\shiftreg_data~56_combout ),
	.datad(address_for_transfer_3),
	.cin(gnd),
	.combout(\shiftreg_data~57_combout ),
	.cout());
defparam \shiftreg_data~57 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~70 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~57_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~70_combout ),
	.cout());
defparam \shiftreg_data~70 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~70 .sum_lutc_input = "datac";

dffeas \shiftreg_data[14] (
	.clk(clk_clk),
	.d(\shiftreg_data~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[14]~q ),
	.prn(vcc));
defparam \shiftreg_data[14] .is_wysiwyg = "true";
defparam \shiftreg_data[14] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~53 (
	.dataa(\shiftreg_data[13]~26_combout ),
	.datab(data_out_15),
	.datac(\shiftreg_data[13]~40_combout ),
	.datad(\shiftreg_data[14]~q ),
	.cin(gnd),
	.combout(\shiftreg_data~53_combout ),
	.cout());
defparam \shiftreg_data~53 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~54 (
	.dataa(address_for_transfer_5),
	.datab(\shiftreg_data[13]~26_combout ),
	.datac(\shiftreg_data~53_combout ),
	.datad(address_for_transfer_4),
	.cin(gnd),
	.combout(\shiftreg_data~54_combout ),
	.cout());
defparam \shiftreg_data~54 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~69 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~54_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~69_combout ),
	.cout());
defparam \shiftreg_data~69 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~69 .sum_lutc_input = "datac";

dffeas \shiftreg_data[15] (
	.clk(clk_clk),
	.d(\shiftreg_data~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[15]~q ),
	.prn(vcc));
defparam \shiftreg_data[15] .is_wysiwyg = "true";
defparam \shiftreg_data[15] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~50 (
	.dataa(\shiftreg_data[13]~40_combout ),
	.datab(address_for_transfer_6),
	.datac(\shiftreg_data[13]~26_combout ),
	.datad(\shiftreg_data[15]~q ),
	.cin(gnd),
	.combout(\shiftreg_data~50_combout ),
	.cout());
defparam \shiftreg_data~50 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~51 (
	.dataa(data_out_16),
	.datab(\shiftreg_data[13]~40_combout ),
	.datac(\shiftreg_data~50_combout ),
	.datad(address_for_transfer_5),
	.cin(gnd),
	.combout(\shiftreg_data~51_combout ),
	.cout());
defparam \shiftreg_data~51 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~68 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~51_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~68_combout ),
	.cout());
defparam \shiftreg_data~68 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~68 .sum_lutc_input = "datac";

dffeas \shiftreg_data[16] (
	.clk(clk_clk),
	.d(\shiftreg_data~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[16]~q ),
	.prn(vcc));
defparam \shiftreg_data[16] .is_wysiwyg = "true";
defparam \shiftreg_data[16] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~47 (
	.dataa(\shiftreg_data[13]~26_combout ),
	.datab(data_out_17),
	.datac(\shiftreg_data[13]~40_combout ),
	.datad(\shiftreg_data[16]~q ),
	.cin(gnd),
	.combout(\shiftreg_data~47_combout ),
	.cout());
defparam \shiftreg_data~47 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~48 (
	.dataa(address_for_transfer_7),
	.datab(\shiftreg_data[13]~26_combout ),
	.datac(\shiftreg_data~47_combout ),
	.datad(address_for_transfer_6),
	.cin(gnd),
	.combout(\shiftreg_data~48_combout ),
	.cout());
defparam \shiftreg_data~48 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~67 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~48_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~67_combout ),
	.cout());
defparam \shiftreg_data~67 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~67 .sum_lutc_input = "datac";

dffeas \shiftreg_data[17] (
	.clk(clk_clk),
	.d(\shiftreg_data~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shiftreg_mask[23]~4_combout ),
	.q(\shiftreg_data[17]~q ),
	.prn(vcc));
defparam \shiftreg_data[17] .is_wysiwyg = "true";
defparam \shiftreg_data[17] .power_up = "low";

cycloneive_lcell_comb \shiftreg_data~23 (
	.dataa(shiftreg_mask),
	.datab(\shiftreg_data[17]~q ),
	.datac(\always4~0_combout ),
	.datad(\s_serial_protocol.STATE_1_INITIALIZE~q ),
	.cin(gnd),
	.combout(\shiftreg_data~23_combout ),
	.cout());
defparam \shiftreg_data~23 .lut_mask = 16'hDFFF;
defparam \shiftreg_data~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~41 (
	.dataa(\shiftreg_data[13]~40_combout ),
	.datab(address_for_transfer_0),
	.datac(\shiftreg_data[13]~26_combout ),
	.datad(shiftreg_data_9),
	.cin(gnd),
	.combout(\shiftreg_data~41_combout ),
	.cout());
defparam \shiftreg_data~41 .lut_mask = 16'hFFDE;
defparam \shiftreg_data~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~42 (
	.dataa(data_out_10),
	.datab(\shiftreg_data[13]~40_combout ),
	.datac(\shiftreg_data~41_combout ),
	.datad(data_reg_8),
	.cin(gnd),
	.combout(\shiftreg_data~42_combout ),
	.cout());
defparam \shiftreg_data~42 .lut_mask = 16'hFFBE;
defparam \shiftreg_data~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \shiftreg_data~66 (
	.dataa(\Serial_Config_Clock_Generator|middle_of_high_level~q ),
	.datab(\s_serial_protocol.STATE_2_RESTART_BIT~q ),
	.datac(shiftreg_mask),
	.datad(\shiftreg_data~42_combout ),
	.cin(gnd),
	.combout(\shiftreg_data~66_combout ),
	.cout());
defparam \shiftreg_data~66 .lut_mask = 16'hFF7F;
defparam \shiftreg_data~66 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_up_slow_clock_generator (
	middle_of_high_level1,
	middle_of_low_level1,
	new_clk1,
	internal_reset,
	internal_reset1,
	r_sync_rst,
	shiftreg_mask,
	clk)/* synthesis synthesis_greybox=1 */;
output 	middle_of_high_level1;
output 	middle_of_low_level1;
output 	new_clk1;
input 	internal_reset;
input 	internal_reset1;
input 	r_sync_rst;
input 	shiftreg_mask;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_counter[1]~11_combout ;
wire \clk_counter[1]~q ;
wire \clk_counter[1]~12 ;
wire \clk_counter[2]~13_combout ;
wire \clk_counter[2]~q ;
wire \clk_counter[2]~14 ;
wire \clk_counter[3]~15_combout ;
wire \clk_counter[3]~q ;
wire \clk_counter[3]~16 ;
wire \clk_counter[4]~17_combout ;
wire \clk_counter[4]~q ;
wire \clk_counter[4]~18 ;
wire \clk_counter[5]~19_combout ;
wire \clk_counter[5]~q ;
wire \clk_counter[5]~20 ;
wire \clk_counter[6]~21_combout ;
wire \clk_counter[6]~q ;
wire \clk_counter[6]~22 ;
wire \clk_counter[7]~23_combout ;
wire \clk_counter[7]~q ;
wire \clk_counter[7]~24 ;
wire \clk_counter[8]~25_combout ;
wire \clk_counter[8]~q ;
wire \clk_counter[8]~26 ;
wire \clk_counter[9]~27_combout ;
wire \clk_counter[9]~q ;
wire \clk_counter[9]~28 ;
wire \clk_counter[10]~29_combout ;
wire \clk_counter[10]~q ;
wire \clk_counter[10]~30 ;
wire \clk_counter[11]~31_combout ;
wire \clk_counter[11]~q ;
wire \middle_of_high_level~0_combout ;
wire \middle_of_high_level~1_combout ;
wire \middle_of_high_level~2_combout ;
wire \middle_of_high_level~3_combout ;
wire \middle_of_low_level~0_combout ;
wire \new_clk~0_combout ;


dffeas middle_of_high_level(
	.clk(clk),
	.d(\middle_of_high_level~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(middle_of_high_level1),
	.prn(vcc));
defparam middle_of_high_level.is_wysiwyg = "true";
defparam middle_of_high_level.power_up = "low";

dffeas middle_of_low_level(
	.clk(clk),
	.d(\middle_of_low_level~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(middle_of_low_level1),
	.prn(vcc));
defparam middle_of_low_level.is_wysiwyg = "true";
defparam middle_of_low_level.power_up = "low";

dffeas new_clk(
	.clk(clk),
	.d(\new_clk~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(new_clk1),
	.prn(vcc));
defparam new_clk.is_wysiwyg = "true";
defparam new_clk.power_up = "low";

cycloneive_lcell_comb \clk_counter[1]~11 (
	.dataa(\clk_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\clk_counter[1]~11_combout ),
	.cout(\clk_counter[1]~12 ));
defparam \clk_counter[1]~11 .lut_mask = 16'h55AA;
defparam \clk_counter[1]~11 .sum_lutc_input = "datac";

dffeas \clk_counter[1] (
	.clk(clk),
	.d(\clk_counter[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[1]~q ),
	.prn(vcc));
defparam \clk_counter[1] .is_wysiwyg = "true";
defparam \clk_counter[1] .power_up = "low";

cycloneive_lcell_comb \clk_counter[2]~13 (
	.dataa(\clk_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[1]~12 ),
	.combout(\clk_counter[2]~13_combout ),
	.cout(\clk_counter[2]~14 ));
defparam \clk_counter[2]~13 .lut_mask = 16'h5A5F;
defparam \clk_counter[2]~13 .sum_lutc_input = "cin";

dffeas \clk_counter[2] (
	.clk(clk),
	.d(\clk_counter[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[2]~q ),
	.prn(vcc));
defparam \clk_counter[2] .is_wysiwyg = "true";
defparam \clk_counter[2] .power_up = "low";

cycloneive_lcell_comb \clk_counter[3]~15 (
	.dataa(\clk_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[2]~14 ),
	.combout(\clk_counter[3]~15_combout ),
	.cout(\clk_counter[3]~16 ));
defparam \clk_counter[3]~15 .lut_mask = 16'h5AAF;
defparam \clk_counter[3]~15 .sum_lutc_input = "cin";

dffeas \clk_counter[3] (
	.clk(clk),
	.d(\clk_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[3]~q ),
	.prn(vcc));
defparam \clk_counter[3] .is_wysiwyg = "true";
defparam \clk_counter[3] .power_up = "low";

cycloneive_lcell_comb \clk_counter[4]~17 (
	.dataa(\clk_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[3]~16 ),
	.combout(\clk_counter[4]~17_combout ),
	.cout(\clk_counter[4]~18 ));
defparam \clk_counter[4]~17 .lut_mask = 16'h5A5F;
defparam \clk_counter[4]~17 .sum_lutc_input = "cin";

dffeas \clk_counter[4] (
	.clk(clk),
	.d(\clk_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[4]~q ),
	.prn(vcc));
defparam \clk_counter[4] .is_wysiwyg = "true";
defparam \clk_counter[4] .power_up = "low";

cycloneive_lcell_comb \clk_counter[5]~19 (
	.dataa(\clk_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[4]~18 ),
	.combout(\clk_counter[5]~19_combout ),
	.cout(\clk_counter[5]~20 ));
defparam \clk_counter[5]~19 .lut_mask = 16'h5AAF;
defparam \clk_counter[5]~19 .sum_lutc_input = "cin";

dffeas \clk_counter[5] (
	.clk(clk),
	.d(\clk_counter[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[5]~q ),
	.prn(vcc));
defparam \clk_counter[5] .is_wysiwyg = "true";
defparam \clk_counter[5] .power_up = "low";

cycloneive_lcell_comb \clk_counter[6]~21 (
	.dataa(\clk_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[5]~20 ),
	.combout(\clk_counter[6]~21_combout ),
	.cout(\clk_counter[6]~22 ));
defparam \clk_counter[6]~21 .lut_mask = 16'h5A5F;
defparam \clk_counter[6]~21 .sum_lutc_input = "cin";

dffeas \clk_counter[6] (
	.clk(clk),
	.d(\clk_counter[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[6]~q ),
	.prn(vcc));
defparam \clk_counter[6] .is_wysiwyg = "true";
defparam \clk_counter[6] .power_up = "low";

cycloneive_lcell_comb \clk_counter[7]~23 (
	.dataa(\clk_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[6]~22 ),
	.combout(\clk_counter[7]~23_combout ),
	.cout(\clk_counter[7]~24 ));
defparam \clk_counter[7]~23 .lut_mask = 16'h5AAF;
defparam \clk_counter[7]~23 .sum_lutc_input = "cin";

dffeas \clk_counter[7] (
	.clk(clk),
	.d(\clk_counter[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[7]~q ),
	.prn(vcc));
defparam \clk_counter[7] .is_wysiwyg = "true";
defparam \clk_counter[7] .power_up = "low";

cycloneive_lcell_comb \clk_counter[8]~25 (
	.dataa(\clk_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[7]~24 ),
	.combout(\clk_counter[8]~25_combout ),
	.cout(\clk_counter[8]~26 ));
defparam \clk_counter[8]~25 .lut_mask = 16'h5A5F;
defparam \clk_counter[8]~25 .sum_lutc_input = "cin";

dffeas \clk_counter[8] (
	.clk(clk),
	.d(\clk_counter[8]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[8]~q ),
	.prn(vcc));
defparam \clk_counter[8] .is_wysiwyg = "true";
defparam \clk_counter[8] .power_up = "low";

cycloneive_lcell_comb \clk_counter[9]~27 (
	.dataa(\clk_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[8]~26 ),
	.combout(\clk_counter[9]~27_combout ),
	.cout(\clk_counter[9]~28 ));
defparam \clk_counter[9]~27 .lut_mask = 16'h5AAF;
defparam \clk_counter[9]~27 .sum_lutc_input = "cin";

dffeas \clk_counter[9] (
	.clk(clk),
	.d(\clk_counter[9]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[9]~q ),
	.prn(vcc));
defparam \clk_counter[9] .is_wysiwyg = "true";
defparam \clk_counter[9] .power_up = "low";

cycloneive_lcell_comb \clk_counter[10]~29 (
	.dataa(\clk_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\clk_counter[9]~28 ),
	.combout(\clk_counter[10]~29_combout ),
	.cout(\clk_counter[10]~30 ));
defparam \clk_counter[10]~29 .lut_mask = 16'h5A5F;
defparam \clk_counter[10]~29 .sum_lutc_input = "cin";

dffeas \clk_counter[10] (
	.clk(clk),
	.d(\clk_counter[10]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[10]~q ),
	.prn(vcc));
defparam \clk_counter[10] .is_wysiwyg = "true";
defparam \clk_counter[10] .power_up = "low";

cycloneive_lcell_comb \clk_counter[11]~31 (
	.dataa(\clk_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\clk_counter[10]~30 ),
	.combout(\clk_counter[11]~31_combout ),
	.cout());
defparam \clk_counter[11]~31 .lut_mask = 16'h5A5A;
defparam \clk_counter[11]~31 .sum_lutc_input = "cin";

dffeas \clk_counter[11] (
	.clk(clk),
	.d(\clk_counter[11]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(shiftreg_mask),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_counter[11]~q ),
	.prn(vcc));
defparam \clk_counter[11] .is_wysiwyg = "true";
defparam \clk_counter[11] .power_up = "low";

cycloneive_lcell_comb \middle_of_high_level~0 (
	.dataa(\clk_counter[3]~q ),
	.datab(\clk_counter[2]~q ),
	.datac(\clk_counter[1]~q ),
	.datad(\clk_counter[10]~q ),
	.cin(gnd),
	.combout(\middle_of_high_level~0_combout ),
	.cout());
defparam \middle_of_high_level~0 .lut_mask = 16'hFEFF;
defparam \middle_of_high_level~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \middle_of_high_level~1 (
	.dataa(\clk_counter[7]~q ),
	.datab(\clk_counter[6]~q ),
	.datac(\clk_counter[5]~q ),
	.datad(\clk_counter[4]~q ),
	.cin(gnd),
	.combout(\middle_of_high_level~1_combout ),
	.cout());
defparam \middle_of_high_level~1 .lut_mask = 16'hFFFE;
defparam \middle_of_high_level~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \middle_of_high_level~2 (
	.dataa(\clk_counter[9]~q ),
	.datab(\clk_counter[8]~q ),
	.datac(\middle_of_high_level~0_combout ),
	.datad(\middle_of_high_level~1_combout ),
	.cin(gnd),
	.combout(\middle_of_high_level~2_combout ),
	.cout());
defparam \middle_of_high_level~2 .lut_mask = 16'hFFFE;
defparam \middle_of_high_level~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \middle_of_high_level~3 (
	.dataa(\clk_counter[11]~q ),
	.datab(\middle_of_high_level~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\middle_of_high_level~3_combout ),
	.cout());
defparam \middle_of_high_level~3 .lut_mask = 16'hEEEE;
defparam \middle_of_high_level~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \middle_of_low_level~0 (
	.dataa(\middle_of_high_level~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\clk_counter[11]~q ),
	.cin(gnd),
	.combout(\middle_of_low_level~0_combout ),
	.cout());
defparam \middle_of_low_level~0 .lut_mask = 16'hAAFF;
defparam \middle_of_low_level~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \new_clk~0 (
	.dataa(\clk_counter[11]~q ),
	.datab(internal_reset),
	.datac(internal_reset1),
	.datad(r_sync_rst),
	.cin(gnd),
	.combout(\new_clk~0_combout ),
	.cout());
defparam \new_clk~0 .lut_mask = 16'hBFFF;
defparam \new_clk~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_audio_pll_0 (
	locked,
	clk_0,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	locked;
output 	clk_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_up_altpll audio_pll(
	.locked(locked),
	.clk_0(clk_0),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_up_altpll (
	locked,
	clk_0,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	locked;
output 	clk_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altpll_1 PLL_for_DE_Series_Boards(
	.locked(locked),
	.clk_0(clk_0),
	.inclk({gnd,clk_clk}));

endmodule

module final_project_soc_altpll_1 (
	locked,
	clk_0,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	locked;
output 	clk_0;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altpll_dkb2 auto_generated(
	.locked(locked),
	.clk({clk_unconnected_wire_5,clk_unconnected_wire_4,clk_unconnected_wire_3,clk_unconnected_wire_2,clk_unconnected_wire_1,clk_0}),
	.inclk({gnd,inclk[0]}));

endmodule

module final_project_soc_altpll_dkb2 (
	locked,
	clk,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	locked;
output 	[5:0] clk;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk[1] ;
wire \clk[2] ;
wire \clk[3] ;
wire \clk[4] ;
wire \pll1~FBOUT ;

wire [4:0] pll1_CLK_bus;

assign clk[0] = pll1_CLK_bus[0];
assign \clk[1]  = pll1_CLK_bus[1];
assign \clk[2]  = pll1_CLK_bus[2];
assign \clk[3]  = pll1_CLK_bus[3];
assign \clk[4]  = pll1_CLK_bus[4];

cycloneive_pll pll1(
	.areset(gnd),
	.pfdena(vcc),
	.fbin(\pll1~FBOUT ),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scandata(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect(3'b000),
	.phasedone(),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(locked),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(\pll1~FBOUT ),
	.clk(pll1_CLK_bus),
	.clkbad());
defparam pll1.auto_settings = "false";
defparam pll1.bandwidth_type = "auto";
defparam pll1.c0_high = 31;
defparam pll1.c0_initial = 1;
defparam pll1.c0_low = 30;
defparam pll1.c0_mode = "odd";
defparam pll1.c0_ph = 0;
defparam pll1.c1_high = 8;
defparam pll1.c1_initial = 1;
defparam pll1.c1_low = 7;
defparam pll1.c1_mode = "odd";
defparam pll1.c1_ph = 0;
defparam pll1.c1_use_casc_in = "off";
defparam pll1.c2_high = 8;
defparam pll1.c2_initial = 1;
defparam pll1.c2_low = 7;
defparam pll1.c2_mode = "odd";
defparam pll1.c2_ph = 0;
defparam pll1.c2_use_casc_in = "off";
defparam pll1.c3_high = 1;
defparam pll1.c3_initial = 1;
defparam pll1.c3_low = 1;
defparam pll1.c3_mode = "bypass";
defparam pll1.c3_ph = 0;
defparam pll1.c3_use_casc_in = "off";
defparam pll1.c4_high = 1;
defparam pll1.c4_initial = 1;
defparam pll1.c4_low = 1;
defparam pll1.c4_mode = "bypass";
defparam pll1.c4_ph = 0;
defparam pll1.c4_use_casc_in = "off";
defparam pll1.charge_pump_current_bits = 2;
defparam pll1.clk0_counter = "c0";
defparam pll1.clk0_divide_by = 297;
defparam pll1.clk0_duty_cycle = 50;
defparam pll1.clk0_multiply_by = 73;
defparam pll1.clk0_phase_shift = "0";
defparam pll1.clk1_counter = "c1";
defparam pll1.clk1_divide_by = 1;
defparam pll1.clk1_duty_cycle = 50;
defparam pll1.clk1_multiply_by = 1;
defparam pll1.clk1_phase_shift = "0";
defparam pll1.clk2_counter = "c2";
defparam pll1.clk2_divide_by = 1;
defparam pll1.clk2_duty_cycle = 50;
defparam pll1.clk2_multiply_by = 1;
defparam pll1.clk2_phase_shift = "0";
defparam pll1.clk3_counter = "unused";
defparam pll1.clk3_divide_by = 0;
defparam pll1.clk3_duty_cycle = 50;
defparam pll1.clk3_multiply_by = 0;
defparam pll1.clk3_phase_shift = "0";
defparam pll1.clk4_counter = "unused";
defparam pll1.clk4_divide_by = 0;
defparam pll1.clk4_duty_cycle = 50;
defparam pll1.clk4_multiply_by = 0;
defparam pll1.clk4_phase_shift = "0";
defparam pll1.compensate_clock = "clock0";
defparam pll1.inclk0_input_frequency = 20000;
defparam pll1.inclk1_input_frequency = 0;
defparam pll1.loop_filter_c_bits = 2;
defparam pll1.loop_filter_r_bits = 1;
defparam pll1.m = 15;
defparam pll1.m_initial = 1;
defparam pll1.m_ph = 0;
defparam pll1.n = 1;
defparam pll1.operation_mode = "normal";
defparam pll1.pfd_max = 0;
defparam pll1.pfd_min = 0;
defparam pll1.self_reset_on_loss_lock = "off";
defparam pll1.simulation_type = "timing";
defparam pll1.switch_over_type = "auto";
defparam pll1.vco_center = 0;
defparam pll1.vco_divide_by = 0;
defparam pll1.vco_frequency_control = "auto";
defparam pll1.vco_max = 0;
defparam pll1.vco_min = 0;
defparam pll1.vco_multiply_by = 0;
defparam pll1.vco_phase_shift_step = 0;
defparam pll1.vco_post_scale = 1;

endmodule

module final_project_soc_final_project_soc_jtag_uart_0 (
	W_alu_result_2,
	tdo,
	d_read,
	d_write,
	read_accepted,
	write_accepted,
	cp_valid,
	uav_write,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	Equal2,
	d_writedata_10,
	uav_read,
	rst1,
	Equal21,
	av_waitrequest1,
	mem_used_1,
	av_readdata_9,
	av_readdata_8,
	b_full,
	read_01,
	av_readdata_0,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_01,
	counter_reg_bit_11,
	counter_reg_bit_41,
	counter_reg_bit_51,
	av_readdata_1,
	av_readdata_2,
	av_readdata_3,
	av_readdata_4,
	av_readdata_5,
	av_readdata_6,
	av_readdata_7,
	ac1,
	woverflow1,
	rvalid1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
output 	tdo;
input 	d_read;
input 	d_write;
input 	read_accepted;
input 	write_accepted;
input 	cp_valid;
input 	uav_write;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	Equal2;
input 	d_writedata_10;
input 	uav_read;
output 	rst1;
input 	Equal21;
output 	av_waitrequest1;
input 	mem_used_1;
output 	av_readdata_9;
output 	av_readdata_8;
output 	b_full;
output 	read_01;
output 	av_readdata_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	counter_reg_bit_31;
output 	counter_reg_bit_21;
output 	counter_reg_bit_01;
output 	counter_reg_bit_11;
output 	counter_reg_bit_41;
output 	counter_reg_bit_51;
output 	av_readdata_1;
output 	av_readdata_2;
output 	av_readdata_3;
output 	av_readdata_4;
output 	av_readdata_5;
output 	av_readdata_6;
output 	av_readdata_7;
output 	ac1;
output 	woverflow1;
output 	rvalid1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ;
wire \t_dav~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_pause~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_ena~q ;
wire \the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_wr~q ;
wire \wr_rfifo~combout ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ;
wire \final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ;
wire \fifo_wr~0_combout ;
wire \av_waitrequest~0_combout ;
wire \av_waitrequest~1_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \ien_AF~2_combout ;
wire \ien_AE~q ;
wire \ien_AF~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~0_combout ;
wire \Add0~2_combout ;
wire \LessThan1~0_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \LessThan1~1_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \LessThan1~2_combout ;
wire \fifo_AF~q ;
wire \fifo_rd~3_combout ;
wire \ac~0_combout ;
wire \ac~1_combout ;
wire \woverflow~3_combout ;
wire \woverflow~2_combout ;
wire \fifo_rd~2_combout ;
wire \rvalid~0_combout ;


final_project_soc_alt_jtag_atlantic final_project_soc_jtag_uart_0_alt_jtag_atlantic(
	.r_dat({\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ,\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ,
\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ,\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ,
\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ,\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ,
\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ,\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] }),
	.tdo1(tdo),
	.rst_n(r_sync_rst),
	.rst11(rst1),
	.t_dav(\t_dav~q ),
	.rvalid01(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.t_pause1(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_pause~q ),
	.t_ena1(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.wdata_0(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

final_project_soc_final_project_soc_jtag_uart_0_scfifo_r the_final_project_soc_jtag_uart_0_scfifo_r(
	.q_b_0(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ),
	.q_b_1(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ),
	.q_b_2(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ),
	.q_b_3(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ),
	.q_b_4(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ),
	.q_b_5(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ),
	.q_b_6(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ),
	.q_b_7(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_31),
	.counter_reg_bit_2(counter_reg_bit_21),
	.counter_reg_bit_0(counter_reg_bit_01),
	.counter_reg_bit_1(counter_reg_bit_11),
	.counter_reg_bit_4(counter_reg_bit_41),
	.counter_reg_bit_5(counter_reg_bit_51),
	.t_ena(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.fifo_rd(\fifo_rd~2_combout ),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_jtag_uart_0_scfifo_w the_final_project_soc_jtag_uart_0_scfifo_w(
	.q_b_7(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ),
	.q_b_0(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ),
	.q_b_1(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ),
	.q_b_2(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ),
	.q_b_3(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ),
	.q_b_4(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ),
	.q_b_5(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ),
	.q_b_6(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.fifo_wr(\fifo_wr~q ),
	.clk_clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

cycloneive_lcell_comb \r_val~0 (
	.dataa(\the_final_project_soc_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datab(\r_val~q ),
	.datac(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.datad(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.cin(gnd),
	.combout(\r_val~0_combout ),
	.cout());
defparam \r_val~0 .lut_mask = 16'hBFFF;
defparam \r_val~0 .sum_lutc_input = "datac";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cycloneive_lcell_comb wr_rfifo(
	.dataa(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(b_full),
	.cin(gnd),
	.combout(\wr_rfifo~combout ),
	.cout());
defparam wr_rfifo.lut_mask = 16'hAAFF;
defparam wr_rfifo.sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_wr~0 (
	.dataa(W_alu_result_2),
	.datab(b_full1),
	.datac(uav_write),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(\fifo_wr~0_combout ),
	.cout());
defparam \fifo_wr~0 .lut_mask = 16'hFFF7;
defparam \fifo_wr~0 .sum_lutc_input = "datac";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

cycloneive_lcell_comb \av_readdata[9] (
	.dataa(\fifo_AE~q ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_9),
	.cout());
defparam \av_readdata[9] .lut_mask = 16'hEEEE;
defparam \av_readdata[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[8]~0 (
	.dataa(\ien_AF~q ),
	.datab(\pause_irq~q ),
	.datac(\fifo_AF~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_8),
	.cout());
defparam \av_readdata[8]~0 .lut_mask = 16'hFEFE;
defparam \av_readdata[8]~0 .sum_lutc_input = "datac";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

cycloneive_lcell_comb \av_readdata[0]~1 (
	.dataa(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[0] ),
	.datab(\ien_AF~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_0),
	.cout());
defparam \av_readdata[0]~1 .lut_mask = 16'hAACC;
defparam \av_readdata[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[1]~2 (
	.dataa(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[1] ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_1),
	.cout());
defparam \av_readdata[1]~2 .lut_mask = 16'hAACC;
defparam \av_readdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[2]~3 (
	.dataa(read_01),
	.datab(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_2),
	.cout());
defparam \av_readdata[2]~3 .lut_mask = 16'hEEEE;
defparam \av_readdata[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[3]~4 (
	.dataa(read_01),
	.datab(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_3),
	.cout());
defparam \av_readdata[3]~4 .lut_mask = 16'hEEEE;
defparam \av_readdata[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[4]~5 (
	.dataa(read_01),
	.datab(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_4),
	.cout());
defparam \av_readdata[4]~5 .lut_mask = 16'hEEEE;
defparam \av_readdata[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[5]~6 (
	.dataa(read_01),
	.datab(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_5),
	.cout());
defparam \av_readdata[5]~6 .lut_mask = 16'hEEEE;
defparam \av_readdata[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[6]~7 (
	.dataa(read_01),
	.datab(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_6),
	.cout());
defparam \av_readdata[6]~7 .lut_mask = 16'hEEEE;
defparam \av_readdata[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[7]~8 (
	.dataa(read_01),
	.datab(\the_final_project_soc_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|altsyncram1|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_7),
	.cout());
defparam \av_readdata[7]~8 .lut_mask = 16'hEEEE;
defparam \av_readdata[7]~8 .sum_lutc_input = "datac";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(Equal2),
	.datab(Equal21),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hEFFF;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~1 (
	.dataa(cp_valid),
	.datab(\av_waitrequest~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest~1_combout ),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'hEEEE;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hFFFE;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\LessThan0~0_combout ),
	.datab(b_full1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cycloneive_lcell_comb \ien_AF~2 (
	.dataa(d_write),
	.datab(write_accepted),
	.datac(W_alu_result_2),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(\ien_AF~2_combout ),
	.cout());
defparam \ien_AF~2 .lut_mask = 16'hFFFB;
defparam \ien_AF~2 .sum_lutc_input = "datac";

dffeas ien_AE(
	.clk(clk_clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~2_combout ),
	.q(\ien_AE~q ),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

dffeas ien_AF(
	.clk(clk_clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~2_combout ),
	.q(\ien_AF~q ),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cycloneive_lcell_comb \pause_irq~0 (
	.dataa(b_non_empty),
	.datab(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_pause~q ),
	.datac(\pause_irq~q ),
	.datad(read_01),
	.cin(gnd),
	.combout(\pause_irq~0_combout ),
	.cout());
defparam \pause_irq~0 .lut_mask = 16'hFEFF;
defparam \pause_irq~0 .sum_lutc_input = "datac";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(counter_reg_bit_01),
	.datab(counter_reg_bit_11),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h6677;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~2 (
	.dataa(counter_reg_bit_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5AAF;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(counter_reg_bit_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5A5F;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~0 (
	.dataa(\Add0~4_combout ),
	.datab(counter_reg_bit_01),
	.datac(\Add0~0_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hFFFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~6 (
	.dataa(counter_reg_bit_41),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5AAF;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~8 (
	.dataa(counter_reg_bit_51),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~1 (
	.dataa(\Add0~6_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
defparam \LessThan1~1 .lut_mask = 16'hEEEE;
defparam \LessThan1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~10 (
	.dataa(b_full),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5AAF;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'hF0F0;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~2 (
	.dataa(\LessThan1~0_combout ),
	.datab(\LessThan1~1_combout ),
	.datac(\Add0~10_combout ),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\LessThan1~2_combout ),
	.cout());
defparam \LessThan1~2 .lut_mask = 16'h7FFF;
defparam \LessThan1~2 .sum_lutc_input = "datac";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cycloneive_lcell_comb \fifo_rd~3 (
	.dataa(d_read),
	.datab(read_accepted),
	.datac(\av_waitrequest~0_combout ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\fifo_rd~3_combout ),
	.cout());
defparam \fifo_rd~3 .lut_mask = 16'hFBFF;
defparam \fifo_rd~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~0 (
	.dataa(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_pause~q ),
	.datab(\final_project_soc_jtag_uart_0_alt_jtag_atlantic|t_ena~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac~0_combout ),
	.cout());
defparam \ac~0 .lut_mask = 16'hEEEE;
defparam \ac~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~1 (
	.dataa(\ac~0_combout ),
	.datab(ac1),
	.datac(d_writedata_10),
	.datad(\ien_AF~2_combout ),
	.cin(gnd),
	.combout(\ac~1_combout ),
	.cout());
defparam \ac~1 .lut_mask = 16'hEFFF;
defparam \ac~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~3 (
	.dataa(d_write),
	.datab(write_accepted),
	.datac(\av_waitrequest~0_combout ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\woverflow~3_combout ),
	.cout());
defparam \woverflow~3 .lut_mask = 16'hFBFF;
defparam \woverflow~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~2 (
	.dataa(b_full1),
	.datab(woverflow1),
	.datac(gnd),
	.datad(\woverflow~3_combout ),
	.cin(gnd),
	.combout(\woverflow~2_combout ),
	.cout());
defparam \woverflow~2 .lut_mask = 16'hAACC;
defparam \woverflow~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_rd~2 (
	.dataa(uav_read),
	.datab(\av_waitrequest~0_combout ),
	.datac(b_non_empty),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\fifo_rd~2_combout ),
	.cout());
defparam \fifo_rd~2 .lut_mask = 16'hFEFF;
defparam \fifo_rd~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rvalid~0 (
	.dataa(\fifo_rd~2_combout ),
	.datab(rvalid1),
	.datac(gnd),
	.datad(\fifo_rd~3_combout ),
	.cin(gnd),
	.combout(\rvalid~0_combout ),
	.cout());
defparam \rvalid~0 .lut_mask = 16'hEEFF;
defparam \rvalid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_alt_jtag_atlantic (
	r_dat,
	tdo1,
	rst_n,
	rst11,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_pause1,
	t_ena1,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	tdo1;
input 	rst_n;
output 	rst11;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_pause1;
output 	t_ena1;
output 	wdata_0;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	wdata_6;
output 	wdata_7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \count~2_combout ;
wire \td_shift[0]~4_combout ;
wire \count[1]~q ;
wire \count~10_combout ;
wire \count[2]~q ;
wire \count~9_combout ;
wire \count[3]~q ;
wire \count~8_combout ;
wire \count[4]~q ;
wire \count~7_combout ;
wire \count[5]~q ;
wire \count~6_combout ;
wire \count[6]~q ;
wire \count~5_combout ;
wire \count[7]~q ;
wire \count~3_combout ;
wire \count[8]~q ;
wire \always0~0_combout ;
wire \state~0_combout ;
wire \state~1_combout ;
wire \state~2_combout ;
wire \state~q ;
wire \count[9]~0_combout ;
wire \count[9]~1_combout ;
wire \count[9]~q ;
wire \count~4_combout ;
wire \count[0]~q ;
wire \wdata[1]~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~1_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift~11_combout ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~8_combout ;
wire \td_shift[9]~q ;
wire \td_shift~6_combout ;
wire \rdata[6]~q ;
wire \td_shift~22_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~20_combout ;
wire \td_shift~21_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~18_combout ;
wire \td_shift~19_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~16_combout ;
wire \td_shift~17_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~14_combout ;
wire \td_shift~15_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~12_combout ;
wire \td_shift~13_combout ;
wire \td_shift[3]~q ;
wire \rdata[0]~q ;
wire \td_shift~9_combout ;
wire \td_shift~10_combout ;
wire \td_shift[2]~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~2_combout ;
wire \write_stalled~q ;
wire \td_shift~5_combout ;
wire \td_shift~7_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~0_combout ;
wire \td_shift~1_combout ;
wire \td_shift~2_combout ;
wire \td_shift~3_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \read_req~q ;
wire \rvalid0~1_combout ;
wire \rst2~q ;
wire \rvalid0~2_combout ;
wire \write~0_combout ;
wire \wdata[1]~1_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~0_combout ;
wire \write_valid~q ;
wire \t_pause~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \t_pause~1_combout ;
wire \t_ena~2_combout ;
wire \t_ena~3_combout ;


dffeas tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tdo1),
	.prn(vcc));
defparam tdo.is_wysiwyg = "true";
defparam tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~2_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas t_pause(
	.clk(clk),
	.d(\t_pause~1_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause1),
	.prn(vcc));
defparam t_pause.is_wysiwyg = "true";
defparam t_pause.power_up = "low";

dffeas t_ena(
	.clk(clk),
	.d(\t_ena~3_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena1),
	.prn(vcc));
defparam t_ena.is_wysiwyg = "true";
defparam t_ena.power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

cycloneive_lcell_comb \tck_t_dav~0 (
	.dataa(t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tck_t_dav~0_combout ),
	.cout());
defparam \tck_t_dav~0 .lut_mask = 16'h5555;
defparam \tck_t_dav~0 .sum_lutc_input = "datac";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cycloneive_lcell_comb \count~2 (
	.dataa(state_4),
	.datab(\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~2_combout ),
	.cout());
defparam \count~2 .lut_mask = 16'hEEEE;
defparam \count~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift[0]~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(state_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\td_shift[0]~4_combout ),
	.cout());
defparam \td_shift[0]~4 .lut_mask = 16'hFEFF;
defparam \td_shift[0]~4 .sum_lutc_input = "datac";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \count~10 (
	.dataa(\count[1]~q ),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~10_combout ),
	.cout());
defparam \count~10 .lut_mask = 16'hEEEE;
defparam \count~10 .sum_lutc_input = "datac";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count~9 (
	.dataa(state_4),
	.datab(\count[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~9_combout ),
	.cout());
defparam \count~9 .lut_mask = 16'hEEEE;
defparam \count~9 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count~8 (
	.dataa(state_4),
	.datab(\count[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~8_combout ),
	.cout());
defparam \count~8 .lut_mask = 16'hEEEE;
defparam \count~8 .sum_lutc_input = "datac";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count~7 (
	.dataa(state_4),
	.datab(\count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~7_combout ),
	.cout());
defparam \count~7 .lut_mask = 16'hEEEE;
defparam \count~7 .sum_lutc_input = "datac";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count~6 (
	.dataa(state_4),
	.datab(\count[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~6_combout ),
	.cout());
defparam \count~6 .lut_mask = 16'hEEEE;
defparam \count~6 .sum_lutc_input = "datac";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count~5 (
	.dataa(state_4),
	.datab(\count[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEEEE;
defparam \count~5 .sum_lutc_input = "datac";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \count~3 (
	.dataa(state_4),
	.datab(\count[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hEEEE;
defparam \count~3 .sum_lutc_input = "datac";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(gnd),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~0 (
	.dataa(state_4),
	.datab(\always0~0_combout ),
	.datac(altera_internal_jtag1),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hFEFF;
defparam \state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~1 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'h7777;
defparam \state~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~2 (
	.dataa(\state~q ),
	.datab(virtual_ir_scan_reg),
	.datac(\state~0_combout ),
	.datad(\state~1_combout ),
	.cin(gnd),
	.combout(\state~2_combout ),
	.cout());
defparam \state~2 .lut_mask = 16'hFFD8;
defparam \state~2 .sum_lutc_input = "datac";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cycloneive_lcell_comb \count[9]~0 (
	.dataa(altera_internal_jtag1),
	.datab(irf_reg_0_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[9]~0_combout ),
	.cout());
defparam \count[9]~0 .lut_mask = 16'hBBBB;
defparam \count[9]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[9]~1 (
	.dataa(state_4),
	.datab(\count[8]~q ),
	.datac(\state~q ),
	.datad(\count[9]~0_combout ),
	.cin(gnd),
	.combout(\count[9]~1_combout ),
	.cout());
defparam \count[9]~1 .lut_mask = 16'hF7FF;
defparam \count[9]~1 .sum_lutc_input = "datac";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cycloneive_lcell_comb \count~4 (
	.dataa(state_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hAAFF;
defparam \count~4 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \wdata[1]~0 (
	.dataa(\state~q ),
	.datab(state_4),
	.datac(splitter_nodes_receive_0_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\wdata[1]~0_combout ),
	.cout());
defparam \wdata[1]~0 .lut_mask = 16'hFEFF;
defparam \wdata[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \user_saw_rvalid~0 (
	.dataa(\td_shift[0]~q ),
	.datab(\user_saw_rvalid~q ),
	.datac(irf_reg_0_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.cout());
defparam \user_saw_rvalid~0 .lut_mask = 16'hACAC;
defparam \user_saw_rvalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \user_saw_rvalid~1 (
	.dataa(\user_saw_rvalid~q ),
	.datab(\count[0]~q ),
	.datac(\wdata[1]~0_combout ),
	.datad(\user_saw_rvalid~0_combout ),
	.cin(gnd),
	.combout(\user_saw_rvalid~1_combout ),
	.cout());
defparam \user_saw_rvalid~1 .lut_mask = 16'hFFBE;
defparam \user_saw_rvalid~1 .sum_lutc_input = "datac";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~11 (
	.dataa(altera_internal_jtag1),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~11_combout ),
	.cout());
defparam \td_shift~11 .lut_mask = 16'hEEEE;
defparam \td_shift~11 .sum_lutc_input = "datac";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cycloneive_lcell_comb \r_ena~0 (
	.dataa(r_val),
	.datab(r_ena11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\r_ena~0_combout ),
	.cout());
defparam \r_ena~0 .lut_mask = 16'hEEEE;
defparam \r_ena~0 .sum_lutc_input = "datac";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cycloneive_lcell_comb \td_shift~8 (
	.dataa(\td_shift[10]~q ),
	.datab(\rdata[7]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~8_combout ),
	.cout());
defparam \td_shift~8 .lut_mask = 16'hAACC;
defparam \td_shift~8 .sum_lutc_input = "datac";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cycloneive_lcell_comb \td_shift~6 (
	.dataa(\user_saw_rvalid~q ),
	.datab(\td_shift[9]~q ),
	.datac(\state~q ),
	.datad(\count[1]~q ),
	.cin(gnd),
	.combout(\td_shift~6_combout ),
	.cout());
defparam \td_shift~6 .lut_mask = 16'hEFFF;
defparam \td_shift~6 .sum_lutc_input = "datac";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cycloneive_lcell_comb \td_shift~22 (
	.dataa(\td_shift[9]~q ),
	.datab(\rdata[6]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~22_combout ),
	.cout());
defparam \td_shift~22 .lut_mask = 16'hAACC;
defparam \td_shift~22 .sum_lutc_input = "datac";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~22_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cycloneive_lcell_comb \td_shift~20 (
	.dataa(\td_shift[8]~q ),
	.datab(\rdata[5]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~20_combout ),
	.cout());
defparam \td_shift~20 .lut_mask = 16'hACAC;
defparam \td_shift~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~21 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(\td_shift~20_combout ),
	.cin(gnd),
	.combout(\td_shift~21_combout ),
	.cout());
defparam \td_shift~21 .lut_mask = 16'hFFFE;
defparam \td_shift~21 .sum_lutc_input = "datac";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~21_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cycloneive_lcell_comb \td_shift~18 (
	.dataa(\td_shift[7]~q ),
	.datab(\rdata[4]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~18_combout ),
	.cout());
defparam \td_shift~18 .lut_mask = 16'hAACC;
defparam \td_shift~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~19 (
	.dataa(\td_shift~18_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~19_combout ),
	.cout());
defparam \td_shift~19 .lut_mask = 16'hFAFC;
defparam \td_shift~19 .sum_lutc_input = "datac";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~19_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cycloneive_lcell_comb \td_shift~16 (
	.dataa(\td_shift[6]~q ),
	.datab(\rdata[3]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~16_combout ),
	.cout());
defparam \td_shift~16 .lut_mask = 16'hAACC;
defparam \td_shift~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~17 (
	.dataa(\td_shift~16_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~17_combout ),
	.cout());
defparam \td_shift~17 .lut_mask = 16'hFAFC;
defparam \td_shift~17 .sum_lutc_input = "datac";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~17_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cycloneive_lcell_comb \td_shift~14 (
	.dataa(\td_shift[5]~q ),
	.datab(\rdata[2]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~14_combout ),
	.cout());
defparam \td_shift~14 .lut_mask = 16'hACAC;
defparam \td_shift~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~15 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(\td_shift~14_combout ),
	.cin(gnd),
	.combout(\td_shift~15_combout ),
	.cout());
defparam \td_shift~15 .lut_mask = 16'hFFFE;
defparam \td_shift~15 .sum_lutc_input = "datac";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~15_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cycloneive_lcell_comb \td_shift~12 (
	.dataa(\td_shift[4]~q ),
	.datab(\rdata[1]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~12_combout ),
	.cout());
defparam \td_shift~12 .lut_mask = 16'hACAC;
defparam \td_shift~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~13 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(\td_shift~12_combout ),
	.cin(gnd),
	.combout(\td_shift~13_combout ),
	.cout());
defparam \td_shift~13 .lut_mask = 16'hFFFE;
defparam \td_shift~13 .sum_lutc_input = "datac";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~13_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

cycloneive_lcell_comb \td_shift~9 (
	.dataa(\td_shift[3]~q ),
	.datab(\rdata[0]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~9_combout ),
	.cout());
defparam \td_shift~9 .lut_mask = 16'hAACC;
defparam \td_shift~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~10 (
	.dataa(\td_shift~9_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~10_combout ),
	.cout());
defparam \td_shift~10 .lut_mask = 16'hFAFC;
defparam \td_shift~10 .sum_lutc_input = "datac";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cycloneive_lcell_comb \write_stalled~0 (
	.dataa(\td_shift[10]~q ),
	.datab(\write_stalled~q ),
	.datac(\tck_t_dav~q ),
	.datad(altera_internal_jtag1),
	.cin(gnd),
	.combout(\write_stalled~0_combout ),
	.cout());
defparam \write_stalled~0 .lut_mask = 16'hEFFF;
defparam \write_stalled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~1 (
	.dataa(state_4),
	.datab(splitter_nodes_receive_0_3),
	.datac(virtual_ir_scan_reg),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_stalled~1_combout ),
	.cout());
defparam \write_stalled~1 .lut_mask = 16'hEFEF;
defparam \write_stalled~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~2 (
	.dataa(\count[1]~q ),
	.datab(irf_reg_0_1),
	.datac(\state~q ),
	.datad(\write_stalled~1_combout ),
	.cin(gnd),
	.combout(\write_stalled~2_combout ),
	.cout());
defparam \write_stalled~2 .lut_mask = 16'hFFFB;
defparam \write_stalled~2 .sum_lutc_input = "datac";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cycloneive_lcell_comb \td_shift~5 (
	.dataa(\td_shift[2]~q ),
	.datab(\write_stalled~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~5_combout ),
	.cout());
defparam \td_shift~5 .lut_mask = 16'hAACC;
defparam \td_shift~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~7 (
	.dataa(\td_shift~5_combout ),
	.datab(irf_reg_0_1),
	.datac(\td_shift~6_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\td_shift~7_combout ),
	.cout());
defparam \td_shift~7 .lut_mask = 16'hFAFC;
defparam \td_shift~7 .sum_lutc_input = "datac";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~0 (
	.dataa(\td_shift[1]~q ),
	.datab(\rvalid~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~0_combout ),
	.cout());
defparam \td_shift~0 .lut_mask = 16'hACAC;
defparam \td_shift~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~1 (
	.dataa(\user_saw_rvalid~q ),
	.datab(\td_shift[9]~q ),
	.datac(\count[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~1_combout ),
	.cout());
defparam \td_shift~1 .lut_mask = 16'hF7F7;
defparam \td_shift~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~2 (
	.dataa(\state~q ),
	.datab(altera_internal_jtag1),
	.datac(irf_reg_0_1),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~2_combout ),
	.cout());
defparam \td_shift~2 .lut_mask = 16'hDF8F;
defparam \td_shift~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~3 (
	.dataa(\tck_t_dav~q ),
	.datab(\td_shift~0_combout ),
	.datac(\state~q ),
	.datad(\td_shift~2_combout ),
	.cin(gnd),
	.combout(\td_shift~3_combout ),
	.cout());
defparam \td_shift~3 .lut_mask = 16'hAFCF;
defparam \td_shift~3 .sum_lutc_input = "datac";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cycloneive_lcell_comb \rvalid0~0 (
	.dataa(rvalid01),
	.datab(r_val),
	.datac(r_ena11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rvalid0~0_combout ),
	.cout());
defparam \rvalid0~0 .lut_mask = 16'h7F7F;
defparam \rvalid0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h5555;
defparam \read~0 .sum_lutc_input = "datac";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cycloneive_lcell_comb \rvalid0~1 (
	.dataa(\read1~q ),
	.datab(\read2~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\read_req~q ),
	.cin(gnd),
	.combout(\rvalid0~1_combout ),
	.cout());
defparam \rvalid0~1 .lut_mask = 16'h6FFF;
defparam \rvalid0~1 .sum_lutc_input = "datac";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cycloneive_lcell_comb \rvalid0~2 (
	.dataa(\rvalid0~0_combout ),
	.datab(\rvalid0~1_combout ),
	.datac(gnd),
	.datad(\rst2~q ),
	.cin(gnd),
	.combout(\rvalid0~2_combout ),
	.cout());
defparam \rvalid0~2 .lut_mask = 16'hDDFF;
defparam \rvalid0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~0 (
	.dataa(\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'h5555;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wdata[1]~1 (
	.dataa(\count[8]~q ),
	.datab(irf_reg_0_1),
	.datac(\state~q ),
	.datad(\write_stalled~1_combout ),
	.cin(gnd),
	.combout(\wdata[1]~1_combout ),
	.cout());
defparam \wdata[1]~1 .lut_mask = 16'hFFFB;
defparam \wdata[1]~1 .sum_lutc_input = "datac";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~1_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cycloneive_lcell_comb \always2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\write1~q ),
	.datad(\write2~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h0FF0;
defparam \always2~0 .sum_lutc_input = "datac";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~2_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cycloneive_lcell_comb \t_pause~0 (
	.dataa(\always2~0_combout ),
	.datab(t_dav),
	.datac(\write_stalled~q ),
	.datad(\write_valid~q ),
	.cin(gnd),
	.combout(\t_pause~0_combout ),
	.cout());
defparam \t_pause~0 .lut_mask = 16'hFEFF;
defparam \t_pause~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jupdate~0 (
	.dataa(\jupdate~q ),
	.datab(irf_reg_0_1),
	.datac(\always0~0_combout ),
	.datad(state_8),
	.cin(gnd),
	.combout(\jupdate~0_combout ),
	.cout());
defparam \jupdate~0 .lut_mask = 16'h6996;
defparam \jupdate~0 .sum_lutc_input = "datac";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cycloneive_lcell_comb \t_pause~1 (
	.dataa(\rst2~q ),
	.datab(\t_pause~0_combout ),
	.datac(\jupdate1~q ),
	.datad(\jupdate2~q ),
	.cin(gnd),
	.combout(\t_pause~1_combout ),
	.cout());
defparam \t_pause~1 .lut_mask = 16'hEFFE;
defparam \t_pause~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_ena~2 (
	.dataa(t_ena1),
	.datab(\write_valid~q ),
	.datac(t_dav),
	.datad(\write_stalled~q ),
	.cin(gnd),
	.combout(\t_ena~2_combout ),
	.cout());
defparam \t_ena~2 .lut_mask = 16'hEFFF;
defparam \t_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_ena~3 (
	.dataa(\write1~q ),
	.datab(\write2~q ),
	.datac(\rst2~q ),
	.datad(\t_ena~2_combout ),
	.cin(gnd),
	.combout(\t_ena~3_combout ),
	.cout());
defparam \t_ena~3 .lut_mask = 16'hFFF6;
defparam \t_ena~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_jtag_uart_0_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	fifo_rd,
	wr_rfifo,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	fifo_rd;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_6;
input 	wdata_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_5 rfifo(
	.q({q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,
q_unconnected_wire_19,q_unconnected_wire_18,q_unconnected_wire_17,q_unconnected_wire_16,q_unconnected_wire_15,q_unconnected_wire_14,q_unconnected_wire_13,q_unconnected_wire_12,q_unconnected_wire_11,q_unconnected_wire_10,q_unconnected_wire_9,q_unconnected_wire_8,q_b_7,
q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wr_rfifo),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module final_project_soc_scfifo_5 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[31:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_jr21 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module final_project_soc_scfifo_jr21 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_a_dpfifo_q131 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module final_project_soc_a_dpfifo_q131 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	fifo_rd,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


final_project_soc_cntr_1ob_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

final_project_soc_cntr_1ob rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

final_project_soc_dpram_nl21 FIFOram(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.outclocken(fifo_rd),
	.wren(wreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wraddress({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.rdaddress({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.outclock(clock));

final_project_soc_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wreq),
	.clock(clock));

endmodule

module final_project_soc_a_fefifo_7cf (
	r_sync_rst,
	b_full1,
	b_non_empty1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	t_ena,
	fifo_rd,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	b_non_empty1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \b_non_empty~1_combout ;


final_project_soc_cntr_do7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_5(counter_reg_bit_5),
	.updown(wreq),
	._(\_~4_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~4 (
	.dataa(t_ena),
	.datab(b_full1),
	.datac(fifo_rd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'h9696;
defparam \_~4 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cycloneive_lcell_comb \b_full~0 (
	.dataa(b_non_empty1),
	.datab(counter_reg_bit_3),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_5),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_1),
	.datad(t_ena),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(fifo_rd),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(b_full1),
	.datab(t_ena),
	.datac(gnd),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hEEFF;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_4),
	.datab(counter_reg_bit_5),
	.datac(wreq),
	.datad(\_~2_combout ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFFFE;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(\b_non_empty~0_combout ),
	.datab(b_non_empty1),
	.datac(\_~3_combout ),
	.datad(fifo_rd),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hFEFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_cntr_do7 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_5,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_1ob (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_1ob_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_dpram_nl21 (
	q,
	outclocken,
	wren,
	data,
	wraddress,
	rdaddress,
	outclock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	outclocken;
input 	wren;
input 	[7:0] data;
input 	[5:0] wraddress;
input 	[5:0] rdaddress;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_r1m1 altsyncram1(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(outclocken),
	.wren_a(wren),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({wraddress[5],wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.address_b({rdaddress[5],rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.clock1(outclock),
	.clock0(outclock));

endmodule

module final_project_soc_altsyncram_r1m1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block2a0_PORTBDATAOUT_bus;
wire [143:0] ram_block2a1_PORTBDATAOUT_bus;
wire [143:0] ram_block2a2_PORTBDATAOUT_bus;
wire [143:0] ram_block2a3_PORTBDATAOUT_bus;
wire [143:0] ram_block2a4_PORTBDATAOUT_bus;
wire [143:0] ram_block2a5_PORTBDATAOUT_bus;
wire [143:0] ram_block2a6_PORTBDATAOUT_bus;
wire [143:0] ram_block2a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block2a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block2a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block2a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block2a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block2a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block2a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block2a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block2a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block2a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a0_PORTBDATAOUT_bus));
defparam ram_block2a0.clk0_core_clock_enable = "ena0";
defparam ram_block2a0.clk1_core_clock_enable = "ena1";
defparam ram_block2a0.clk1_input_clock_enable = "ena1";
defparam ram_block2a0.data_interleave_offset_in_bits = 1;
defparam ram_block2a0.data_interleave_width_in_bits = 1;
defparam ram_block2a0.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a0.operation_mode = "dual_port";
defparam ram_block2a0.port_a_address_clear = "none";
defparam ram_block2a0.port_a_address_width = 6;
defparam ram_block2a0.port_a_data_out_clear = "none";
defparam ram_block2a0.port_a_data_out_clock = "none";
defparam ram_block2a0.port_a_data_width = 1;
defparam ram_block2a0.port_a_first_address = 0;
defparam ram_block2a0.port_a_first_bit_number = 0;
defparam ram_block2a0.port_a_last_address = 63;
defparam ram_block2a0.port_a_logical_ram_depth = 64;
defparam ram_block2a0.port_a_logical_ram_width = 8;
defparam ram_block2a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_address_clear = "none";
defparam ram_block2a0.port_b_address_clock = "clock1";
defparam ram_block2a0.port_b_address_width = 6;
defparam ram_block2a0.port_b_data_out_clear = "none";
defparam ram_block2a0.port_b_data_out_clock = "none";
defparam ram_block2a0.port_b_data_width = 1;
defparam ram_block2a0.port_b_first_address = 0;
defparam ram_block2a0.port_b_first_bit_number = 0;
defparam ram_block2a0.port_b_last_address = 63;
defparam ram_block2a0.port_b_logical_ram_depth = 64;
defparam ram_block2a0.port_b_logical_ram_width = 8;
defparam ram_block2a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_read_enable_clock = "clock1";
defparam ram_block2a0.ram_block_type = "auto";

cycloneive_ram_block ram_block2a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a1_PORTBDATAOUT_bus));
defparam ram_block2a1.clk0_core_clock_enable = "ena0";
defparam ram_block2a1.clk1_core_clock_enable = "ena1";
defparam ram_block2a1.clk1_input_clock_enable = "ena1";
defparam ram_block2a1.data_interleave_offset_in_bits = 1;
defparam ram_block2a1.data_interleave_width_in_bits = 1;
defparam ram_block2a1.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a1.operation_mode = "dual_port";
defparam ram_block2a1.port_a_address_clear = "none";
defparam ram_block2a1.port_a_address_width = 6;
defparam ram_block2a1.port_a_data_out_clear = "none";
defparam ram_block2a1.port_a_data_out_clock = "none";
defparam ram_block2a1.port_a_data_width = 1;
defparam ram_block2a1.port_a_first_address = 0;
defparam ram_block2a1.port_a_first_bit_number = 1;
defparam ram_block2a1.port_a_last_address = 63;
defparam ram_block2a1.port_a_logical_ram_depth = 64;
defparam ram_block2a1.port_a_logical_ram_width = 8;
defparam ram_block2a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_address_clear = "none";
defparam ram_block2a1.port_b_address_clock = "clock1";
defparam ram_block2a1.port_b_address_width = 6;
defparam ram_block2a1.port_b_data_out_clear = "none";
defparam ram_block2a1.port_b_data_out_clock = "none";
defparam ram_block2a1.port_b_data_width = 1;
defparam ram_block2a1.port_b_first_address = 0;
defparam ram_block2a1.port_b_first_bit_number = 1;
defparam ram_block2a1.port_b_last_address = 63;
defparam ram_block2a1.port_b_logical_ram_depth = 64;
defparam ram_block2a1.port_b_logical_ram_width = 8;
defparam ram_block2a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_read_enable_clock = "clock1";
defparam ram_block2a1.ram_block_type = "auto";

cycloneive_ram_block ram_block2a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a2_PORTBDATAOUT_bus));
defparam ram_block2a2.clk0_core_clock_enable = "ena0";
defparam ram_block2a2.clk1_core_clock_enable = "ena1";
defparam ram_block2a2.clk1_input_clock_enable = "ena1";
defparam ram_block2a2.data_interleave_offset_in_bits = 1;
defparam ram_block2a2.data_interleave_width_in_bits = 1;
defparam ram_block2a2.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a2.operation_mode = "dual_port";
defparam ram_block2a2.port_a_address_clear = "none";
defparam ram_block2a2.port_a_address_width = 6;
defparam ram_block2a2.port_a_data_out_clear = "none";
defparam ram_block2a2.port_a_data_out_clock = "none";
defparam ram_block2a2.port_a_data_width = 1;
defparam ram_block2a2.port_a_first_address = 0;
defparam ram_block2a2.port_a_first_bit_number = 2;
defparam ram_block2a2.port_a_last_address = 63;
defparam ram_block2a2.port_a_logical_ram_depth = 64;
defparam ram_block2a2.port_a_logical_ram_width = 8;
defparam ram_block2a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_address_clear = "none";
defparam ram_block2a2.port_b_address_clock = "clock1";
defparam ram_block2a2.port_b_address_width = 6;
defparam ram_block2a2.port_b_data_out_clear = "none";
defparam ram_block2a2.port_b_data_out_clock = "none";
defparam ram_block2a2.port_b_data_width = 1;
defparam ram_block2a2.port_b_first_address = 0;
defparam ram_block2a2.port_b_first_bit_number = 2;
defparam ram_block2a2.port_b_last_address = 63;
defparam ram_block2a2.port_b_logical_ram_depth = 64;
defparam ram_block2a2.port_b_logical_ram_width = 8;
defparam ram_block2a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_read_enable_clock = "clock1";
defparam ram_block2a2.ram_block_type = "auto";

cycloneive_ram_block ram_block2a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a3_PORTBDATAOUT_bus));
defparam ram_block2a3.clk0_core_clock_enable = "ena0";
defparam ram_block2a3.clk1_core_clock_enable = "ena1";
defparam ram_block2a3.clk1_input_clock_enable = "ena1";
defparam ram_block2a3.data_interleave_offset_in_bits = 1;
defparam ram_block2a3.data_interleave_width_in_bits = 1;
defparam ram_block2a3.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a3.operation_mode = "dual_port";
defparam ram_block2a3.port_a_address_clear = "none";
defparam ram_block2a3.port_a_address_width = 6;
defparam ram_block2a3.port_a_data_out_clear = "none";
defparam ram_block2a3.port_a_data_out_clock = "none";
defparam ram_block2a3.port_a_data_width = 1;
defparam ram_block2a3.port_a_first_address = 0;
defparam ram_block2a3.port_a_first_bit_number = 3;
defparam ram_block2a3.port_a_last_address = 63;
defparam ram_block2a3.port_a_logical_ram_depth = 64;
defparam ram_block2a3.port_a_logical_ram_width = 8;
defparam ram_block2a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_address_clear = "none";
defparam ram_block2a3.port_b_address_clock = "clock1";
defparam ram_block2a3.port_b_address_width = 6;
defparam ram_block2a3.port_b_data_out_clear = "none";
defparam ram_block2a3.port_b_data_out_clock = "none";
defparam ram_block2a3.port_b_data_width = 1;
defparam ram_block2a3.port_b_first_address = 0;
defparam ram_block2a3.port_b_first_bit_number = 3;
defparam ram_block2a3.port_b_last_address = 63;
defparam ram_block2a3.port_b_logical_ram_depth = 64;
defparam ram_block2a3.port_b_logical_ram_width = 8;
defparam ram_block2a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_read_enable_clock = "clock1";
defparam ram_block2a3.ram_block_type = "auto";

cycloneive_ram_block ram_block2a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a4_PORTBDATAOUT_bus));
defparam ram_block2a4.clk0_core_clock_enable = "ena0";
defparam ram_block2a4.clk1_core_clock_enable = "ena1";
defparam ram_block2a4.clk1_input_clock_enable = "ena1";
defparam ram_block2a4.data_interleave_offset_in_bits = 1;
defparam ram_block2a4.data_interleave_width_in_bits = 1;
defparam ram_block2a4.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a4.operation_mode = "dual_port";
defparam ram_block2a4.port_a_address_clear = "none";
defparam ram_block2a4.port_a_address_width = 6;
defparam ram_block2a4.port_a_data_out_clear = "none";
defparam ram_block2a4.port_a_data_out_clock = "none";
defparam ram_block2a4.port_a_data_width = 1;
defparam ram_block2a4.port_a_first_address = 0;
defparam ram_block2a4.port_a_first_bit_number = 4;
defparam ram_block2a4.port_a_last_address = 63;
defparam ram_block2a4.port_a_logical_ram_depth = 64;
defparam ram_block2a4.port_a_logical_ram_width = 8;
defparam ram_block2a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_address_clear = "none";
defparam ram_block2a4.port_b_address_clock = "clock1";
defparam ram_block2a4.port_b_address_width = 6;
defparam ram_block2a4.port_b_data_out_clear = "none";
defparam ram_block2a4.port_b_data_out_clock = "none";
defparam ram_block2a4.port_b_data_width = 1;
defparam ram_block2a4.port_b_first_address = 0;
defparam ram_block2a4.port_b_first_bit_number = 4;
defparam ram_block2a4.port_b_last_address = 63;
defparam ram_block2a4.port_b_logical_ram_depth = 64;
defparam ram_block2a4.port_b_logical_ram_width = 8;
defparam ram_block2a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_read_enable_clock = "clock1";
defparam ram_block2a4.ram_block_type = "auto";

cycloneive_ram_block ram_block2a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a5_PORTBDATAOUT_bus));
defparam ram_block2a5.clk0_core_clock_enable = "ena0";
defparam ram_block2a5.clk1_core_clock_enable = "ena1";
defparam ram_block2a5.clk1_input_clock_enable = "ena1";
defparam ram_block2a5.data_interleave_offset_in_bits = 1;
defparam ram_block2a5.data_interleave_width_in_bits = 1;
defparam ram_block2a5.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a5.operation_mode = "dual_port";
defparam ram_block2a5.port_a_address_clear = "none";
defparam ram_block2a5.port_a_address_width = 6;
defparam ram_block2a5.port_a_data_out_clear = "none";
defparam ram_block2a5.port_a_data_out_clock = "none";
defparam ram_block2a5.port_a_data_width = 1;
defparam ram_block2a5.port_a_first_address = 0;
defparam ram_block2a5.port_a_first_bit_number = 5;
defparam ram_block2a5.port_a_last_address = 63;
defparam ram_block2a5.port_a_logical_ram_depth = 64;
defparam ram_block2a5.port_a_logical_ram_width = 8;
defparam ram_block2a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_address_clear = "none";
defparam ram_block2a5.port_b_address_clock = "clock1";
defparam ram_block2a5.port_b_address_width = 6;
defparam ram_block2a5.port_b_data_out_clear = "none";
defparam ram_block2a5.port_b_data_out_clock = "none";
defparam ram_block2a5.port_b_data_width = 1;
defparam ram_block2a5.port_b_first_address = 0;
defparam ram_block2a5.port_b_first_bit_number = 5;
defparam ram_block2a5.port_b_last_address = 63;
defparam ram_block2a5.port_b_logical_ram_depth = 64;
defparam ram_block2a5.port_b_logical_ram_width = 8;
defparam ram_block2a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_read_enable_clock = "clock1";
defparam ram_block2a5.ram_block_type = "auto";

cycloneive_ram_block ram_block2a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a6_PORTBDATAOUT_bus));
defparam ram_block2a6.clk0_core_clock_enable = "ena0";
defparam ram_block2a6.clk1_core_clock_enable = "ena1";
defparam ram_block2a6.clk1_input_clock_enable = "ena1";
defparam ram_block2a6.data_interleave_offset_in_bits = 1;
defparam ram_block2a6.data_interleave_width_in_bits = 1;
defparam ram_block2a6.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a6.operation_mode = "dual_port";
defparam ram_block2a6.port_a_address_clear = "none";
defparam ram_block2a6.port_a_address_width = 6;
defparam ram_block2a6.port_a_data_out_clear = "none";
defparam ram_block2a6.port_a_data_out_clock = "none";
defparam ram_block2a6.port_a_data_width = 1;
defparam ram_block2a6.port_a_first_address = 0;
defparam ram_block2a6.port_a_first_bit_number = 6;
defparam ram_block2a6.port_a_last_address = 63;
defparam ram_block2a6.port_a_logical_ram_depth = 64;
defparam ram_block2a6.port_a_logical_ram_width = 8;
defparam ram_block2a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_address_clear = "none";
defparam ram_block2a6.port_b_address_clock = "clock1";
defparam ram_block2a6.port_b_address_width = 6;
defparam ram_block2a6.port_b_data_out_clear = "none";
defparam ram_block2a6.port_b_data_out_clock = "none";
defparam ram_block2a6.port_b_data_width = 1;
defparam ram_block2a6.port_b_first_address = 0;
defparam ram_block2a6.port_b_first_bit_number = 6;
defparam ram_block2a6.port_b_last_address = 63;
defparam ram_block2a6.port_b_logical_ram_depth = 64;
defparam ram_block2a6.port_b_logical_ram_width = 8;
defparam ram_block2a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_read_enable_clock = "clock1";
defparam ram_block2a6.ram_block_type = "auto";

cycloneive_ram_block ram_block2a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a7_PORTBDATAOUT_bus));
defparam ram_block2a7.clk0_core_clock_enable = "ena0";
defparam ram_block2a7.clk1_core_clock_enable = "ena1";
defparam ram_block2a7.clk1_input_clock_enable = "ena1";
defparam ram_block2a7.data_interleave_offset_in_bits = 1;
defparam ram_block2a7.data_interleave_width_in_bits = 1;
defparam ram_block2a7.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_r:the_final_project_soc_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a7.operation_mode = "dual_port";
defparam ram_block2a7.port_a_address_clear = "none";
defparam ram_block2a7.port_a_address_width = 6;
defparam ram_block2a7.port_a_data_out_clear = "none";
defparam ram_block2a7.port_a_data_out_clock = "none";
defparam ram_block2a7.port_a_data_width = 1;
defparam ram_block2a7.port_a_first_address = 0;
defparam ram_block2a7.port_a_first_bit_number = 7;
defparam ram_block2a7.port_a_last_address = 63;
defparam ram_block2a7.port_a_logical_ram_depth = 64;
defparam ram_block2a7.port_a_logical_ram_width = 8;
defparam ram_block2a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_address_clear = "none";
defparam ram_block2a7.port_b_address_clock = "clock1";
defparam ram_block2a7.port_b_address_width = 6;
defparam ram_block2a7.port_b_data_out_clear = "none";
defparam ram_block2a7.port_b_data_out_clock = "none";
defparam ram_block2a7.port_b_data_width = 1;
defparam ram_block2a7.port_b_first_address = 0;
defparam ram_block2a7.port_b_first_bit_number = 7;
defparam ram_block2a7.port_b_last_address = 63;
defparam ram_block2a7.port_b_logical_ram_depth = 64;
defparam ram_block2a7.port_b_logical_ram_width = 8;
defparam ram_block2a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_read_enable_clock = "clock1";
defparam ram_block2a7.ram_block_type = "auto";

endmodule

module final_project_soc_final_project_soc_jtag_uart_0_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	fifo_wr,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	fifo_wr;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_6 wfifo(
	.q({q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,
q_unconnected_wire_19,q_unconnected_wire_18,q_unconnected_wire_17,q_unconnected_wire_16,q_unconnected_wire_15,q_unconnected_wire_14,q_unconnected_wire_13,q_unconnected_wire_12,q_unconnected_wire_11,q_unconnected_wire_10,q_unconnected_wire_9,q_unconnected_wire_8,q_b_7,
q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(fifo_wr),
	.clock(clk_clk));

endmodule

module final_project_soc_scfifo_6 (
	q,
	data,
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	wrreq,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q;
input 	[31:0] data;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_scfifo_jr21_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(wrreq),
	.clock(clock));

endmodule

module final_project_soc_scfifo_jr21_1 (
	q,
	data,
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	wrreq,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_a_dpfifo_q131_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wreq(wrreq),
	.clock(clock));

endmodule

module final_project_soc_a_dpfifo_q131_1 (
	q,
	data,
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	r_val,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
input 	r_val;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


final_project_soc_cntr_1ob_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

final_project_soc_cntr_1ob_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

final_project_soc_dpram_nl21_1 FIFOram(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.outclocken(r_val),
	.wren(wreq),
	.wraddress({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.rdaddress({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.outclock(clock));

final_project_soc_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full1(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.wreq(wreq),
	.clock(clock));

endmodule

module final_project_soc_a_fefifo_7cf_1 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty1,
	r_val,
	wreq,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty1;
input 	r_val;
input 	wreq;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;


final_project_soc_cntr_do7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.updown(wreq),
	._(\_~0_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(wreq),
	.datad(r_val),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FF0;
defparam \_~0 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cycloneive_lcell_comb \b_full~0 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(wreq),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hFFFE;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(counter_reg_bit_3),
	.datab(\b_non_empty~0_combout ),
	.datac(counter_reg_bit_0),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hEFFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~2 (
	.dataa(b_full1),
	.datab(wreq),
	.datac(b_non_empty1),
	.datad(\b_non_empty~1_combout ),
	.cin(gnd),
	.combout(\b_non_empty~2_combout ),
	.cout());
defparam \b_non_empty~2 .lut_mask = 16'hFFFE;
defparam \b_non_empty~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_cntr_do7_1 (
	r_sync_rst,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_1ob_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_cntr_1ob_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module final_project_soc_dpram_nl21_1 (
	q,
	data,
	outclocken,
	wren,
	wraddress,
	rdaddress,
	outclock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	outclocken;
input 	wren;
input 	[5:0] wraddress;
input 	[5:0] rdaddress;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_r1m1_1 altsyncram1(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clocken1(outclocken),
	.wren_a(wren),
	.address_a({wraddress[5],wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.address_b({rdaddress[5],rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.clock1(outclock),
	.clock0(outclock));

endmodule

module final_project_soc_altsyncram_r1m1_1 (
	q_b,
	data_a,
	clocken1,
	wren_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	clocken1;
input 	wren_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block2a7_PORTBDATAOUT_bus;
wire [143:0] ram_block2a0_PORTBDATAOUT_bus;
wire [143:0] ram_block2a1_PORTBDATAOUT_bus;
wire [143:0] ram_block2a2_PORTBDATAOUT_bus;
wire [143:0] ram_block2a3_PORTBDATAOUT_bus;
wire [143:0] ram_block2a4_PORTBDATAOUT_bus;
wire [143:0] ram_block2a5_PORTBDATAOUT_bus;
wire [143:0] ram_block2a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block2a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block2a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block2a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block2a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block2a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block2a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block2a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block2a6_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block2a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a7_PORTBDATAOUT_bus));
defparam ram_block2a7.clk0_core_clock_enable = "ena0";
defparam ram_block2a7.clk1_core_clock_enable = "ena1";
defparam ram_block2a7.clk1_input_clock_enable = "ena1";
defparam ram_block2a7.data_interleave_offset_in_bits = 1;
defparam ram_block2a7.data_interleave_width_in_bits = 1;
defparam ram_block2a7.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a7.operation_mode = "dual_port";
defparam ram_block2a7.port_a_address_clear = "none";
defparam ram_block2a7.port_a_address_width = 6;
defparam ram_block2a7.port_a_data_out_clear = "none";
defparam ram_block2a7.port_a_data_out_clock = "none";
defparam ram_block2a7.port_a_data_width = 1;
defparam ram_block2a7.port_a_first_address = 0;
defparam ram_block2a7.port_a_first_bit_number = 7;
defparam ram_block2a7.port_a_last_address = 63;
defparam ram_block2a7.port_a_logical_ram_depth = 64;
defparam ram_block2a7.port_a_logical_ram_width = 8;
defparam ram_block2a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_address_clear = "none";
defparam ram_block2a7.port_b_address_clock = "clock1";
defparam ram_block2a7.port_b_address_width = 6;
defparam ram_block2a7.port_b_data_out_clear = "none";
defparam ram_block2a7.port_b_data_out_clock = "none";
defparam ram_block2a7.port_b_data_width = 1;
defparam ram_block2a7.port_b_first_address = 0;
defparam ram_block2a7.port_b_first_bit_number = 7;
defparam ram_block2a7.port_b_last_address = 63;
defparam ram_block2a7.port_b_logical_ram_depth = 64;
defparam ram_block2a7.port_b_logical_ram_width = 8;
defparam ram_block2a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a7.port_b_read_enable_clock = "clock1";
defparam ram_block2a7.ram_block_type = "auto";

cycloneive_ram_block ram_block2a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a0_PORTBDATAOUT_bus));
defparam ram_block2a0.clk0_core_clock_enable = "ena0";
defparam ram_block2a0.clk1_core_clock_enable = "ena1";
defparam ram_block2a0.clk1_input_clock_enable = "ena1";
defparam ram_block2a0.data_interleave_offset_in_bits = 1;
defparam ram_block2a0.data_interleave_width_in_bits = 1;
defparam ram_block2a0.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a0.operation_mode = "dual_port";
defparam ram_block2a0.port_a_address_clear = "none";
defparam ram_block2a0.port_a_address_width = 6;
defparam ram_block2a0.port_a_data_out_clear = "none";
defparam ram_block2a0.port_a_data_out_clock = "none";
defparam ram_block2a0.port_a_data_width = 1;
defparam ram_block2a0.port_a_first_address = 0;
defparam ram_block2a0.port_a_first_bit_number = 0;
defparam ram_block2a0.port_a_last_address = 63;
defparam ram_block2a0.port_a_logical_ram_depth = 64;
defparam ram_block2a0.port_a_logical_ram_width = 8;
defparam ram_block2a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_address_clear = "none";
defparam ram_block2a0.port_b_address_clock = "clock1";
defparam ram_block2a0.port_b_address_width = 6;
defparam ram_block2a0.port_b_data_out_clear = "none";
defparam ram_block2a0.port_b_data_out_clock = "none";
defparam ram_block2a0.port_b_data_width = 1;
defparam ram_block2a0.port_b_first_address = 0;
defparam ram_block2a0.port_b_first_bit_number = 0;
defparam ram_block2a0.port_b_last_address = 63;
defparam ram_block2a0.port_b_logical_ram_depth = 64;
defparam ram_block2a0.port_b_logical_ram_width = 8;
defparam ram_block2a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a0.port_b_read_enable_clock = "clock1";
defparam ram_block2a0.ram_block_type = "auto";

cycloneive_ram_block ram_block2a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a1_PORTBDATAOUT_bus));
defparam ram_block2a1.clk0_core_clock_enable = "ena0";
defparam ram_block2a1.clk1_core_clock_enable = "ena1";
defparam ram_block2a1.clk1_input_clock_enable = "ena1";
defparam ram_block2a1.data_interleave_offset_in_bits = 1;
defparam ram_block2a1.data_interleave_width_in_bits = 1;
defparam ram_block2a1.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a1.operation_mode = "dual_port";
defparam ram_block2a1.port_a_address_clear = "none";
defparam ram_block2a1.port_a_address_width = 6;
defparam ram_block2a1.port_a_data_out_clear = "none";
defparam ram_block2a1.port_a_data_out_clock = "none";
defparam ram_block2a1.port_a_data_width = 1;
defparam ram_block2a1.port_a_first_address = 0;
defparam ram_block2a1.port_a_first_bit_number = 1;
defparam ram_block2a1.port_a_last_address = 63;
defparam ram_block2a1.port_a_logical_ram_depth = 64;
defparam ram_block2a1.port_a_logical_ram_width = 8;
defparam ram_block2a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_address_clear = "none";
defparam ram_block2a1.port_b_address_clock = "clock1";
defparam ram_block2a1.port_b_address_width = 6;
defparam ram_block2a1.port_b_data_out_clear = "none";
defparam ram_block2a1.port_b_data_out_clock = "none";
defparam ram_block2a1.port_b_data_width = 1;
defparam ram_block2a1.port_b_first_address = 0;
defparam ram_block2a1.port_b_first_bit_number = 1;
defparam ram_block2a1.port_b_last_address = 63;
defparam ram_block2a1.port_b_logical_ram_depth = 64;
defparam ram_block2a1.port_b_logical_ram_width = 8;
defparam ram_block2a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a1.port_b_read_enable_clock = "clock1";
defparam ram_block2a1.ram_block_type = "auto";

cycloneive_ram_block ram_block2a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a2_PORTBDATAOUT_bus));
defparam ram_block2a2.clk0_core_clock_enable = "ena0";
defparam ram_block2a2.clk1_core_clock_enable = "ena1";
defparam ram_block2a2.clk1_input_clock_enable = "ena1";
defparam ram_block2a2.data_interleave_offset_in_bits = 1;
defparam ram_block2a2.data_interleave_width_in_bits = 1;
defparam ram_block2a2.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a2.operation_mode = "dual_port";
defparam ram_block2a2.port_a_address_clear = "none";
defparam ram_block2a2.port_a_address_width = 6;
defparam ram_block2a2.port_a_data_out_clear = "none";
defparam ram_block2a2.port_a_data_out_clock = "none";
defparam ram_block2a2.port_a_data_width = 1;
defparam ram_block2a2.port_a_first_address = 0;
defparam ram_block2a2.port_a_first_bit_number = 2;
defparam ram_block2a2.port_a_last_address = 63;
defparam ram_block2a2.port_a_logical_ram_depth = 64;
defparam ram_block2a2.port_a_logical_ram_width = 8;
defparam ram_block2a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_address_clear = "none";
defparam ram_block2a2.port_b_address_clock = "clock1";
defparam ram_block2a2.port_b_address_width = 6;
defparam ram_block2a2.port_b_data_out_clear = "none";
defparam ram_block2a2.port_b_data_out_clock = "none";
defparam ram_block2a2.port_b_data_width = 1;
defparam ram_block2a2.port_b_first_address = 0;
defparam ram_block2a2.port_b_first_bit_number = 2;
defparam ram_block2a2.port_b_last_address = 63;
defparam ram_block2a2.port_b_logical_ram_depth = 64;
defparam ram_block2a2.port_b_logical_ram_width = 8;
defparam ram_block2a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a2.port_b_read_enable_clock = "clock1";
defparam ram_block2a2.ram_block_type = "auto";

cycloneive_ram_block ram_block2a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a3_PORTBDATAOUT_bus));
defparam ram_block2a3.clk0_core_clock_enable = "ena0";
defparam ram_block2a3.clk1_core_clock_enable = "ena1";
defparam ram_block2a3.clk1_input_clock_enable = "ena1";
defparam ram_block2a3.data_interleave_offset_in_bits = 1;
defparam ram_block2a3.data_interleave_width_in_bits = 1;
defparam ram_block2a3.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a3.operation_mode = "dual_port";
defparam ram_block2a3.port_a_address_clear = "none";
defparam ram_block2a3.port_a_address_width = 6;
defparam ram_block2a3.port_a_data_out_clear = "none";
defparam ram_block2a3.port_a_data_out_clock = "none";
defparam ram_block2a3.port_a_data_width = 1;
defparam ram_block2a3.port_a_first_address = 0;
defparam ram_block2a3.port_a_first_bit_number = 3;
defparam ram_block2a3.port_a_last_address = 63;
defparam ram_block2a3.port_a_logical_ram_depth = 64;
defparam ram_block2a3.port_a_logical_ram_width = 8;
defparam ram_block2a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_address_clear = "none";
defparam ram_block2a3.port_b_address_clock = "clock1";
defparam ram_block2a3.port_b_address_width = 6;
defparam ram_block2a3.port_b_data_out_clear = "none";
defparam ram_block2a3.port_b_data_out_clock = "none";
defparam ram_block2a3.port_b_data_width = 1;
defparam ram_block2a3.port_b_first_address = 0;
defparam ram_block2a3.port_b_first_bit_number = 3;
defparam ram_block2a3.port_b_last_address = 63;
defparam ram_block2a3.port_b_logical_ram_depth = 64;
defparam ram_block2a3.port_b_logical_ram_width = 8;
defparam ram_block2a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a3.port_b_read_enable_clock = "clock1";
defparam ram_block2a3.ram_block_type = "auto";

cycloneive_ram_block ram_block2a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a4_PORTBDATAOUT_bus));
defparam ram_block2a4.clk0_core_clock_enable = "ena0";
defparam ram_block2a4.clk1_core_clock_enable = "ena1";
defparam ram_block2a4.clk1_input_clock_enable = "ena1";
defparam ram_block2a4.data_interleave_offset_in_bits = 1;
defparam ram_block2a4.data_interleave_width_in_bits = 1;
defparam ram_block2a4.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a4.operation_mode = "dual_port";
defparam ram_block2a4.port_a_address_clear = "none";
defparam ram_block2a4.port_a_address_width = 6;
defparam ram_block2a4.port_a_data_out_clear = "none";
defparam ram_block2a4.port_a_data_out_clock = "none";
defparam ram_block2a4.port_a_data_width = 1;
defparam ram_block2a4.port_a_first_address = 0;
defparam ram_block2a4.port_a_first_bit_number = 4;
defparam ram_block2a4.port_a_last_address = 63;
defparam ram_block2a4.port_a_logical_ram_depth = 64;
defparam ram_block2a4.port_a_logical_ram_width = 8;
defparam ram_block2a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_address_clear = "none";
defparam ram_block2a4.port_b_address_clock = "clock1";
defparam ram_block2a4.port_b_address_width = 6;
defparam ram_block2a4.port_b_data_out_clear = "none";
defparam ram_block2a4.port_b_data_out_clock = "none";
defparam ram_block2a4.port_b_data_width = 1;
defparam ram_block2a4.port_b_first_address = 0;
defparam ram_block2a4.port_b_first_bit_number = 4;
defparam ram_block2a4.port_b_last_address = 63;
defparam ram_block2a4.port_b_logical_ram_depth = 64;
defparam ram_block2a4.port_b_logical_ram_width = 8;
defparam ram_block2a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a4.port_b_read_enable_clock = "clock1";
defparam ram_block2a4.ram_block_type = "auto";

cycloneive_ram_block ram_block2a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a5_PORTBDATAOUT_bus));
defparam ram_block2a5.clk0_core_clock_enable = "ena0";
defparam ram_block2a5.clk1_core_clock_enable = "ena1";
defparam ram_block2a5.clk1_input_clock_enable = "ena1";
defparam ram_block2a5.data_interleave_offset_in_bits = 1;
defparam ram_block2a5.data_interleave_width_in_bits = 1;
defparam ram_block2a5.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a5.operation_mode = "dual_port";
defparam ram_block2a5.port_a_address_clear = "none";
defparam ram_block2a5.port_a_address_width = 6;
defparam ram_block2a5.port_a_data_out_clear = "none";
defparam ram_block2a5.port_a_data_out_clock = "none";
defparam ram_block2a5.port_a_data_width = 1;
defparam ram_block2a5.port_a_first_address = 0;
defparam ram_block2a5.port_a_first_bit_number = 5;
defparam ram_block2a5.port_a_last_address = 63;
defparam ram_block2a5.port_a_logical_ram_depth = 64;
defparam ram_block2a5.port_a_logical_ram_width = 8;
defparam ram_block2a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_address_clear = "none";
defparam ram_block2a5.port_b_address_clock = "clock1";
defparam ram_block2a5.port_b_address_width = 6;
defparam ram_block2a5.port_b_data_out_clear = "none";
defparam ram_block2a5.port_b_data_out_clock = "none";
defparam ram_block2a5.port_b_data_width = 1;
defparam ram_block2a5.port_b_first_address = 0;
defparam ram_block2a5.port_b_first_bit_number = 5;
defparam ram_block2a5.port_b_last_address = 63;
defparam ram_block2a5.port_b_logical_ram_depth = 64;
defparam ram_block2a5.port_b_logical_ram_width = 8;
defparam ram_block2a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a5.port_b_read_enable_clock = "clock1";
defparam ram_block2a5.ram_block_type = "auto";

cycloneive_ram_block ram_block2a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block2a6_PORTBDATAOUT_bus));
defparam ram_block2a6.clk0_core_clock_enable = "ena0";
defparam ram_block2a6.clk1_core_clock_enable = "ena1";
defparam ram_block2a6.clk1_input_clock_enable = "ena1";
defparam ram_block2a6.data_interleave_offset_in_bits = 1;
defparam ram_block2a6.data_interleave_width_in_bits = 1;
defparam ram_block2a6.logical_ram_name = "final_project_soc_jtag_uart_0:jtag_uart_0|final_project_soc_jtag_uart_0_scfifo_w:the_final_project_soc_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_q131:dpfifo|dpram_nl21:FIFOram|altsyncram_r1m1:altsyncram1|ALTSYNCRAM";
defparam ram_block2a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block2a6.operation_mode = "dual_port";
defparam ram_block2a6.port_a_address_clear = "none";
defparam ram_block2a6.port_a_address_width = 6;
defparam ram_block2a6.port_a_data_out_clear = "none";
defparam ram_block2a6.port_a_data_out_clock = "none";
defparam ram_block2a6.port_a_data_width = 1;
defparam ram_block2a6.port_a_first_address = 0;
defparam ram_block2a6.port_a_first_bit_number = 6;
defparam ram_block2a6.port_a_last_address = 63;
defparam ram_block2a6.port_a_logical_ram_depth = 64;
defparam ram_block2a6.port_a_logical_ram_width = 8;
defparam ram_block2a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_address_clear = "none";
defparam ram_block2a6.port_b_address_clock = "clock1";
defparam ram_block2a6.port_b_address_width = 6;
defparam ram_block2a6.port_b_data_out_clear = "none";
defparam ram_block2a6.port_b_data_out_clock = "none";
defparam ram_block2a6.port_b_data_width = 1;
defparam ram_block2a6.port_b_first_address = 0;
defparam ram_block2a6.port_b_first_bit_number = 6;
defparam ram_block2a6.port_b_last_address = 63;
defparam ram_block2a6.port_b_logical_ram_depth = 64;
defparam ram_block2a6.port_b_logical_ram_width = 8;
defparam ram_block2a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block2a6.port_b_read_enable_clock = "clock1";
defparam ram_block2a6.ram_block_type = "auto";

endmodule

module final_project_soc_final_project_soc_LEDG (
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	d_write,
	write_accepted,
	writedata,
	reset_n,
	Equal0,
	mem_used_1,
	always0,
	always01,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	d_write;
input 	write_accepted;
input 	[31:0] writedata;
input 	reset_n;
input 	Equal0;
input 	mem_used_1;
output 	always0;
output 	always01;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~2_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(W_alu_result_7),
	.datab(Equal0),
	.datac(W_alu_result_5),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hEFFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~1 (
	.dataa(d_write),
	.datab(write_accepted),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(always01),
	.cout());
defparam \always0~1 .lut_mask = 16'hBFFF;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAFFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAFFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAFFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAFFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAFFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAFFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAFFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAFFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~2 (
	.dataa(always0),
	.datab(always01),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hEFFF;
defparam \always0~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_LEDR (
	W_alu_result_6,
	W_alu_result_2,
	W_alu_result_3,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	writedata,
	reset_n,
	always0,
	Equal2,
	mem_used_1,
	always01,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_6;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_16;
output 	data_out_17;
input 	[31:0] writedata;
input 	reset_n;
input 	always0;
input 	Equal2;
input 	mem_used_1;
output 	always01;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(writedata[16]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(writedata[17]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(W_alu_result_6),
	.datab(Equal2),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(always01),
	.cout());
defparam \always0~0 .lut_mask = 16'hEEFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAFFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAFFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAFFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAFFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAFFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAFFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAFFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAFFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[8] (
	.dataa(data_out_8),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_8),
	.cout());
defparam \readdata[8] .lut_mask = 16'hAFFF;
defparam \readdata[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[9] (
	.dataa(data_out_9),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_9),
	.cout());
defparam \readdata[9] .lut_mask = 16'hAFFF;
defparam \readdata[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[10] (
	.dataa(data_out_10),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_10),
	.cout());
defparam \readdata[10] .lut_mask = 16'hAFFF;
defparam \readdata[10] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[11] (
	.dataa(data_out_11),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_11),
	.cout());
defparam \readdata[11] .lut_mask = 16'hAFFF;
defparam \readdata[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[12] (
	.dataa(data_out_12),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_12),
	.cout());
defparam \readdata[12] .lut_mask = 16'hAFFF;
defparam \readdata[12] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[13] (
	.dataa(data_out_13),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_13),
	.cout());
defparam \readdata[13] .lut_mask = 16'hAFFF;
defparam \readdata[13] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[14] (
	.dataa(data_out_14),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_14),
	.cout());
defparam \readdata[14] .lut_mask = 16'hAFFF;
defparam \readdata[14] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[15] (
	.dataa(data_out_15),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_15),
	.cout());
defparam \readdata[15] .lut_mask = 16'hAFFF;
defparam \readdata[15] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[16] (
	.dataa(data_out_16),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_16),
	.cout());
defparam \readdata[16] .lut_mask = 16'hAFFF;
defparam \readdata[16] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[17] (
	.dataa(data_out_17),
	.datab(gnd),
	.datac(W_alu_result_2),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(readdata_17),
	.cout());
defparam \readdata[17] .lut_mask = 16'hAFFF;
defparam \readdata[17] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~1 (
	.dataa(always0),
	.datab(always01),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hEFFF;
defparam \always0~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0 (
	wire_pll7_clk_0,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_11,
	W_alu_result_2,
	W_alu_result_3,
	clk_0,
	q_a_0,
	readdata_0,
	q_a_1,
	readdata_1,
	readdata_2,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	readdata_16,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	readdata_17,
	q_a_17,
	q_a_10,
	q_a_9,
	q_a_23,
	readdata_8,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	readdata_01,
	readdata_11,
	readdata_21,
	readdata_3,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	readdata_02,
	readdata_12,
	readdata_22,
	readdata_31,
	readdata_4,
	readdata_111,
	readdata_13,
	readdata_161,
	readdata_121,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_211,
	readdata_18,
	readdata_171,
	readdata_311,
	readdata_30,
	readdata_29,
	readdata_28,
	readdata_27,
	readdata_26,
	readdata_25,
	readdata_10,
	readdata_24,
	readdata_9,
	readdata_23,
	readdata_81,
	readdata_221,
	readdata_7,
	readdata_6,
	readdata_20,
	readdata_19,
	saved_grant_1,
	d_read,
	d_write,
	read_accepted,
	write_accepted,
	cp_valid,
	src_valid,
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_3,
	i_read,
	F_pc_2,
	F_pc_4,
	F_pc_9,
	src1_valid,
	saved_grant_0,
	uav_write,
	mem_used_1,
	internal_reset,
	d_writedata_0,
	d_byteenable_0,
	src_data_32,
	F_pc_0,
	src_data_38,
	F_pc_1,
	src_data_39,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	Equal0,
	mem_used_11,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	Equal2,
	mem_used_12,
	always01,
	wait_latency_counter_11,
	wait_latency_counter_01,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	entries_1,
	entries_0,
	altera_reset_synchronizer_int_chain_out1,
	WideOr1,
	uav_read,
	src_data_68,
	waitrequest,
	Equal21,
	s_serial_transferSTATE_1_PRE_WRITE,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	mem_86_0,
	mem_68_0,
	src0_valid,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	src0_valid1,
	src0_valid2,
	read_latency_shift_reg_04,
	mem_86_01,
	mem_68_01,
	src0_valid3,
	src0_valid4,
	WideOr11,
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	mem_67_04,
	mem_67_05,
	mem_67_06,
	out_data_buffer_67,
	out_data_buffer_671,
	mem_67_07,
	src_payload,
	rst1,
	Equal22,
	av_waitrequest,
	mem_used_13,
	waitrequest1,
	mem_used_14,
	mem_used_15,
	saved_grant_01,
	mem_used_16,
	waitrequest2,
	nios2_qsys_0_data_master_waitrequest,
	src1_valid1,
	src1_valid2,
	src1_valid3,
	src_payload1,
	src_payload2,
	out_valid2,
	out_valid3,
	av_readdatavalid,
	saved_grant_02,
	out_data_buffer_3,
	src_data_381,
	src_data_391,
	WideOr12,
	mem_used_17,
	last_cycle,
	nonposted_write_endofpacket,
	WideOr13,
	src_data_382,
	mem,
	src_data_392,
	last_cycle1,
	saved_grant_11,
	WideOr14,
	src_payload3,
	src_data_681,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	src_data_61,
	src_data_60,
	src_data_383,
	src_data_393,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	out_data_buffer_32,
	out_data_buffer_321,
	out_data_buffer_33,
	out_data_buffer_331,
	out_data_buffer_34,
	out_data_buffer_341,
	out_data_buffer_35,
	out_data_buffer_351,
	m0_read,
	WideOr15,
	local_read,
	mem1,
	WideOr16,
	hbreak_enabled,
	av_readdata_pre_30,
	src_payload4,
	av_readdata_pre_0,
	av_readdata_pre_01,
	out_data_buffer_0,
	out_data_buffer_01,
	av_readdata_pre_1,
	out_data_buffer_1,
	av_readdata_pre_11,
	out_data_buffer_11,
	av_readdata_pre_2,
	out_data_buffer_2,
	out_data_buffer_21,
	av_readdata_pre_3,
	readdata_32,
	out_data_buffer_31,
	out_data_buffer_36,
	av_readdata_pre_4,
	readdata_41,
	out_data_buffer_4,
	out_data_buffer_41,
	src_payload5,
	src_data_682,
	src_payload6,
	d_byteenable_2,
	src_payload7,
	mem2,
	src_data_461,
	av_readdata_pre_111,
	out_data_buffer_111,
	out_data_buffer_112,
	av_readdata_pre_13,
	out_data_buffer_13,
	out_data_buffer_131,
	src_payload8,
	av_readdata_pre_16,
	out_data_buffer_16,
	out_data_buffer_161,
	av_readdata_pre_12,
	out_data_buffer_12,
	out_data_buffer_121,
	readdata_51,
	src_payload9,
	av_readdata_pre_5,
	out_data_buffer_5,
	out_data_buffer_51,
	out_data_buffer_14,
	av_readdata_pre_14,
	out_data_buffer_141,
	av_readdata_pre_15,
	out_data_buffer_15,
	out_data_buffer_151,
	av_readdata_pre_21,
	out_data_buffer_211,
	out_data_buffer_212,
	out_data_buffer_18,
	av_readdata_pre_18,
	out_data_buffer_181,
	av_readdata_pre_17,
	out_data_buffer_17,
	out_data_buffer_171,
	av_readdata_pre_31,
	out_data_buffer_311,
	out_data_buffer_312,
	out_data_buffer_30,
	av_readdata_pre_301,
	out_data_buffer_301,
	av_readdata_pre_29,
	out_data_buffer_29,
	out_data_buffer_291,
	out_data_buffer_28,
	av_readdata_pre_28,
	out_data_buffer_281,
	av_readdata_pre_27,
	out_data_buffer_27,
	out_data_buffer_271,
	out_data_buffer_26,
	av_readdata_pre_26,
	out_data_buffer_261,
	av_readdata_pre_25,
	out_data_buffer_25,
	out_data_buffer_251,
	out_data_buffer_10,
	av_readdata_pre_10,
	out_data_buffer_101,
	out_data_buffer_24,
	av_readdata_pre_24,
	out_data_buffer_241,
	av_readdata_pre_9,
	out_data_buffer_9,
	out_data_buffer_91,
	av_readdata_pre_23,
	out_data_buffer_23,
	out_data_buffer_231,
	out_data_buffer_8,
	av_readdata_pre_8,
	out_data_buffer_81,
	out_data_buffer_22,
	av_readdata_pre_22,
	out_data_buffer_221,
	readdata_71,
	out_data_buffer_7,
	av_readdata_pre_7,
	out_data_buffer_71,
	readdata_61,
	av_readdata_pre_6,
	out_data_buffer_6,
	out_data_buffer_61,
	av_readdata_pre_20,
	out_data_buffer_20,
	out_data_buffer_201,
	av_readdata_pre_19,
	out_data_buffer_19,
	out_data_buffer_191,
	src_payload10,
	src_data_0,
	av_readdata_9,
	av_readdata_8,
	src_payload11,
	src_data_384,
	src_data_394,
	src_data_321,
	readdata_03,
	src_payload12,
	readdata_110,
	src_payload13,
	src_payload14,
	readdata_42,
	src_payload15,
	src_payload16,
	src_data_1,
	src_data_11,
	src_data_2,
	src_data_21,
	src_data_3,
	src_data_31,
	src_data_4,
	src_data_410,
	src_data_5,
	src_data_6,
	src_data_63,
	src_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_111,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	d_byteenable_1,
	d_byteenable_3,
	b_full,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	readdata_112,
	src_payload49,
	src_data_33,
	readdata_131,
	src_payload50,
	src_payload51,
	src_data_34,
	readdata_162,
	src_payload52,
	readdata_122,
	src_payload53,
	readdata_52,
	src_payload54,
	readdata_141,
	readdata_151,
	src_payload55,
	out_data_buffer_282,
	out_data_buffer_283,
	readdata_212,
	d_writedata_21,
	src_payload56,
	d_writedata_18,
	src_payload57,
	readdata_181,
	out_data_buffer_272,
	out_data_buffer_273,
	readdata_172,
	src_payload58,
	src_payload59,
	src_data_35,
	readdata_312,
	out_data_buffer_262,
	out_data_buffer_263,
	src_payload60,
	readdata_301,
	out_data_buffer_252,
	out_data_buffer_253,
	src_payload61,
	readdata_291,
	out_data_buffer_242,
	out_data_buffer_243,
	src_payload62,
	readdata_281,
	src_data_23,
	src_payload63,
	readdata_271,
	src_data_22,
	src_payload64,
	readdata_261,
	src_data_211,
	src_payload65,
	readdata_251,
	src_data_20,
	src_payload66,
	readdata_101,
	src_payload67,
	readdata_241,
	src_data_19,
	src_payload68,
	readdata_91,
	d_writedata_23,
	src_payload69,
	readdata_231,
	src_data_18,
	src_payload70,
	readdata_82,
	d_writedata_22,
	src_payload71,
	readdata_222,
	src_payload72,
	readdata_72,
	src_payload73,
	readdata_62,
	readdata_201,
	d_writedata_20,
	src_payload74,
	readdata_191,
	d_writedata_19,
	src_payload75,
	readdata_04,
	read_0,
	av_readdata_0,
	readdata_05,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_01,
	counter_reg_bit_11,
	counter_reg_bit_41,
	counter_reg_bit_51,
	src_payload76,
	readdata_113,
	av_readdata_1,
	readdata_114,
	readdata_210,
	av_readdata_2,
	readdata_213,
	readdata_33,
	av_readdata_3,
	readdata_34,
	readdata_43,
	av_readdata_4,
	readdata_44,
	readdata_53,
	av_readdata_5,
	readdata_54,
	readdata_63,
	av_readdata_6,
	readdata_64,
	readdata_73,
	av_readdata_7,
	readdata_74,
	readdata_83,
	readdata_92,
	readdata_102,
	ac,
	readdata_115,
	readdata_123,
	readdata_132,
	readdata_142,
	woverflow,
	readdata_152,
	rvalid,
	readdata_163,
	readdata_173,
	src_payload77,
	src_payload78,
	src_data_385,
	src_data_395,
	src_data_401,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_322,
	out_data_buffer_313,
	out_data_buffer_314,
	out_data_buffer_302,
	out_data_buffer_303,
	out_data_buffer_292,
	out_data_buffer_293,
	src_payload79,
	src_payload80,
	src_payload81,
	za_valid,
	out_data_buffer_02,
	out_data_buffer_110,
	src_payload82,
	out_data_buffer_210,
	src_payload83,
	src_payload84,
	src_payload85,
	src_data_331,
	src_payload86,
	src_payload87,
	src_data_341,
	src_payload88,
	src_payload89,
	src_payload90,
	src_payload91,
	src_payload92,
	src_payload93,
	src_payload94,
	src_payload95,
	src_data_351,
	src_payload96,
	src_payload97,
	src_payload98,
	src_payload99,
	src_payload100,
	src_payload101,
	src_payload102,
	src_payload103,
	src_payload104,
	src_payload105,
	src_payload106,
	src_payload107,
	src_payload108,
	src_payload109,
	src_payload110,
	src_payload111,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	src_payload112,
	za_data_11,
	za_data_13,
	za_data_16,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_21,
	za_data_18,
	za_data_17,
	za_data_31,
	za_data_30,
	za_data_29,
	za_data_28,
	za_data_27,
	za_data_26,
	za_data_25,
	za_data_10,
	za_data_24,
	za_data_9,
	za_data_23,
	za_data_8,
	za_data_22,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_19,
	src_payload113,
	src_payload114,
	src_payload115,
	src_payload116,
	src_payload117,
	src_payload118,
	src_payload119,
	src_payload120,
	src_payload121,
	src_payload122,
	src_payload123,
	src_payload124,
	src_payload125,
	src_payload126,
	src_payload127,
	src_payload128,
	src_payload129,
	src_payload130,
	src_payload131,
	src_payload132,
	src_payload133,
	src_payload134,
	src_payload135,
	src_payload136,
	src_payload137,
	src_payload138,
	av_ld_getting_data,
	m0_write,
	src_data_510,
	src_data_71,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_28;
input 	W_alu_result_27;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_24;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_12;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_11;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	clk_0;
input 	q_a_0;
input 	readdata_0;
input 	q_a_1;
input 	readdata_1;
input 	readdata_2;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_11;
input 	q_a_13;
input 	readdata_16;
input 	q_a_16;
input 	q_a_12;
input 	q_a_5;
input 	q_a_14;
input 	q_a_15;
input 	q_a_21;
input 	q_a_18;
input 	readdata_17;
input 	q_a_17;
input 	q_a_10;
input 	q_a_9;
input 	q_a_23;
input 	readdata_8;
input 	q_a_8;
input 	q_a_22;
input 	q_a_7;
input 	q_a_6;
input 	q_a_20;
input 	q_a_19;
input 	readdata_01;
input 	readdata_11;
input 	readdata_21;
input 	readdata_3;
input 	d_writedata_31;
input 	d_writedata_30;
input 	d_writedata_29;
input 	d_writedata_28;
input 	d_writedata_27;
input 	d_writedata_26;
input 	d_writedata_25;
input 	d_writedata_24;
input 	readdata_02;
input 	readdata_12;
input 	readdata_22;
input 	readdata_31;
input 	readdata_4;
input 	readdata_111;
input 	readdata_13;
input 	readdata_161;
input 	readdata_121;
input 	readdata_5;
input 	readdata_14;
input 	readdata_15;
input 	readdata_211;
input 	readdata_18;
input 	readdata_171;
input 	readdata_311;
input 	readdata_30;
input 	readdata_29;
input 	readdata_28;
input 	readdata_27;
input 	readdata_26;
input 	readdata_25;
input 	readdata_10;
input 	readdata_24;
input 	readdata_9;
input 	readdata_23;
input 	readdata_81;
input 	readdata_221;
input 	readdata_7;
input 	readdata_6;
input 	readdata_20;
input 	readdata_19;
output 	saved_grant_1;
input 	d_read;
input 	d_write;
output 	read_accepted;
output 	write_accepted;
output 	cp_valid;
output 	src_valid;
input 	F_pc_26;
input 	F_pc_25;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_3;
input 	i_read;
input 	F_pc_2;
input 	F_pc_4;
input 	F_pc_9;
output 	src1_valid;
output 	saved_grant_0;
output 	uav_write;
output 	mem_used_1;
input 	internal_reset;
input 	d_writedata_0;
input 	d_byteenable_0;
output 	src_data_32;
input 	F_pc_0;
output 	src_data_38;
input 	F_pc_1;
output 	src_data_39;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	Equal0;
output 	mem_used_11;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	Equal2;
output 	mem_used_12;
input 	always01;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	entries_1;
input 	entries_0;
input 	altera_reset_synchronizer_int_chain_out1;
output 	WideOr1;
output 	uav_read;
output 	src_data_68;
input 	waitrequest;
input 	Equal21;
input 	s_serial_transferSTATE_1_PRE_WRITE;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg_01;
output 	mem_86_0;
output 	mem_68_0;
output 	src0_valid;
output 	out_valid;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid1;
output 	read_latency_shift_reg_02;
output 	read_latency_shift_reg_03;
output 	src0_valid1;
output 	src0_valid2;
output 	read_latency_shift_reg_04;
output 	mem_86_01;
output 	mem_68_01;
output 	src0_valid3;
output 	src0_valid4;
output 	WideOr11;
output 	mem_67_0;
output 	mem_67_01;
output 	mem_67_02;
output 	mem_67_03;
output 	mem_67_04;
output 	mem_67_05;
output 	mem_67_06;
output 	out_data_buffer_67;
output 	out_data_buffer_671;
output 	mem_67_07;
output 	src_payload;
input 	rst1;
output 	Equal22;
input 	av_waitrequest;
output 	mem_used_13;
input 	waitrequest1;
output 	mem_used_14;
output 	mem_used_15;
output 	saved_grant_01;
output 	mem_used_16;
input 	waitrequest2;
output 	nios2_qsys_0_data_master_waitrequest;
output 	src1_valid1;
output 	src1_valid2;
output 	src1_valid3;
output 	src_payload1;
output 	src_payload2;
output 	out_valid2;
output 	out_valid3;
output 	av_readdatavalid;
output 	saved_grant_02;
output 	out_data_buffer_3;
output 	src_data_381;
output 	src_data_391;
output 	WideOr12;
output 	mem_used_17;
output 	last_cycle;
output 	nonposted_write_endofpacket;
output 	WideOr13;
output 	src_data_382;
output 	mem;
output 	src_data_392;
output 	last_cycle1;
output 	saved_grant_11;
output 	WideOr14;
output 	src_payload3;
output 	src_data_681;
output 	src_data_48;
output 	src_data_62;
output 	src_data_49;
output 	src_data_51;
output 	src_data_50;
output 	src_data_53;
output 	src_data_52;
output 	src_data_55;
output 	src_data_54;
output 	src_data_57;
output 	src_data_56;
output 	src_data_59;
output 	src_data_58;
output 	src_data_61;
output 	src_data_60;
output 	src_data_383;
output 	src_data_393;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	out_data_buffer_32;
output 	out_data_buffer_321;
output 	out_data_buffer_33;
output 	out_data_buffer_331;
output 	out_data_buffer_34;
output 	out_data_buffer_341;
output 	out_data_buffer_35;
output 	out_data_buffer_351;
output 	m0_read;
output 	WideOr15;
output 	local_read;
output 	mem1;
output 	WideOr16;
input 	hbreak_enabled;
output 	av_readdata_pre_30;
output 	src_payload4;
output 	av_readdata_pre_0;
output 	av_readdata_pre_01;
output 	out_data_buffer_0;
output 	out_data_buffer_01;
output 	av_readdata_pre_1;
output 	out_data_buffer_1;
output 	av_readdata_pre_11;
output 	out_data_buffer_11;
output 	av_readdata_pre_2;
output 	out_data_buffer_2;
output 	out_data_buffer_21;
output 	av_readdata_pre_3;
input 	readdata_32;
output 	out_data_buffer_31;
output 	out_data_buffer_36;
output 	av_readdata_pre_4;
input 	readdata_41;
output 	out_data_buffer_4;
output 	out_data_buffer_41;
output 	src_payload5;
output 	src_data_682;
output 	src_payload6;
input 	d_byteenable_2;
output 	src_payload7;
output 	mem2;
output 	src_data_461;
output 	av_readdata_pre_111;
output 	out_data_buffer_111;
output 	out_data_buffer_112;
output 	av_readdata_pre_13;
output 	out_data_buffer_13;
output 	out_data_buffer_131;
output 	src_payload8;
output 	av_readdata_pre_16;
output 	out_data_buffer_16;
output 	out_data_buffer_161;
output 	av_readdata_pre_12;
output 	out_data_buffer_12;
output 	out_data_buffer_121;
input 	readdata_51;
output 	src_payload9;
output 	av_readdata_pre_5;
output 	out_data_buffer_5;
output 	out_data_buffer_51;
output 	out_data_buffer_14;
output 	av_readdata_pre_14;
output 	out_data_buffer_141;
output 	av_readdata_pre_15;
output 	out_data_buffer_15;
output 	out_data_buffer_151;
output 	av_readdata_pre_21;
output 	out_data_buffer_211;
output 	out_data_buffer_212;
output 	out_data_buffer_18;
output 	av_readdata_pre_18;
output 	out_data_buffer_181;
output 	av_readdata_pre_17;
output 	out_data_buffer_17;
output 	out_data_buffer_171;
output 	av_readdata_pre_31;
output 	out_data_buffer_311;
output 	out_data_buffer_312;
output 	out_data_buffer_30;
output 	av_readdata_pre_301;
output 	out_data_buffer_301;
output 	av_readdata_pre_29;
output 	out_data_buffer_29;
output 	out_data_buffer_291;
output 	out_data_buffer_28;
output 	av_readdata_pre_28;
output 	out_data_buffer_281;
output 	av_readdata_pre_27;
output 	out_data_buffer_27;
output 	out_data_buffer_271;
output 	out_data_buffer_26;
output 	av_readdata_pre_26;
output 	out_data_buffer_261;
output 	av_readdata_pre_25;
output 	out_data_buffer_25;
output 	out_data_buffer_251;
output 	out_data_buffer_10;
output 	av_readdata_pre_10;
output 	out_data_buffer_101;
output 	out_data_buffer_24;
output 	av_readdata_pre_24;
output 	out_data_buffer_241;
output 	av_readdata_pre_9;
output 	out_data_buffer_9;
output 	out_data_buffer_91;
output 	av_readdata_pre_23;
output 	out_data_buffer_23;
output 	out_data_buffer_231;
output 	out_data_buffer_8;
output 	av_readdata_pre_8;
output 	out_data_buffer_81;
output 	out_data_buffer_22;
output 	av_readdata_pre_22;
output 	out_data_buffer_221;
input 	readdata_71;
output 	out_data_buffer_7;
output 	av_readdata_pre_7;
output 	out_data_buffer_71;
input 	readdata_61;
output 	av_readdata_pre_6;
output 	out_data_buffer_6;
output 	out_data_buffer_61;
output 	av_readdata_pre_20;
output 	out_data_buffer_20;
output 	out_data_buffer_201;
output 	av_readdata_pre_19;
output 	out_data_buffer_19;
output 	out_data_buffer_191;
output 	src_payload10;
output 	src_data_0;
input 	av_readdata_9;
input 	av_readdata_8;
output 	src_payload11;
output 	src_data_384;
output 	src_data_394;
output 	src_data_321;
input 	readdata_03;
output 	src_payload12;
input 	readdata_110;
output 	src_payload13;
output 	src_payload14;
input 	readdata_42;
output 	src_payload15;
output 	src_payload16;
output 	src_data_1;
output 	src_data_11;
output 	src_data_2;
output 	src_data_21;
output 	src_data_3;
output 	src_data_31;
output 	src_data_4;
output 	src_data_410;
output 	src_data_5;
output 	src_data_6;
output 	src_data_63;
output 	src_data_7;
output 	src_data_8;
output 	src_data_9;
output 	src_data_10;
output 	src_data_111;
output 	src_data_12;
output 	src_data_13;
output 	src_data_14;
output 	src_data_15;
output 	src_data_16;
output 	src_data_17;
input 	d_byteenable_1;
input 	d_byteenable_3;
input 	b_full;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
output 	src_payload35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	src_payload46;
output 	src_payload47;
output 	src_payload48;
input 	readdata_112;
output 	src_payload49;
output 	src_data_33;
input 	readdata_131;
output 	src_payload50;
output 	src_payload51;
output 	src_data_34;
input 	readdata_162;
output 	src_payload52;
input 	readdata_122;
output 	src_payload53;
input 	readdata_52;
output 	src_payload54;
input 	readdata_141;
input 	readdata_151;
output 	src_payload55;
output 	out_data_buffer_282;
output 	out_data_buffer_283;
input 	readdata_212;
input 	d_writedata_21;
output 	src_payload56;
input 	d_writedata_18;
output 	src_payload57;
input 	readdata_181;
output 	out_data_buffer_272;
output 	out_data_buffer_273;
input 	readdata_172;
output 	src_payload58;
output 	src_payload59;
output 	src_data_35;
input 	readdata_312;
output 	out_data_buffer_262;
output 	out_data_buffer_263;
output 	src_payload60;
input 	readdata_301;
output 	out_data_buffer_252;
output 	out_data_buffer_253;
output 	src_payload61;
input 	readdata_291;
output 	out_data_buffer_242;
output 	out_data_buffer_243;
output 	src_payload62;
input 	readdata_281;
output 	src_data_23;
output 	src_payload63;
input 	readdata_271;
output 	src_data_22;
output 	src_payload64;
input 	readdata_261;
output 	src_data_211;
output 	src_payload65;
input 	readdata_251;
output 	src_data_20;
output 	src_payload66;
input 	readdata_101;
output 	src_payload67;
input 	readdata_241;
output 	src_data_19;
output 	src_payload68;
input 	readdata_91;
input 	d_writedata_23;
output 	src_payload69;
input 	readdata_231;
output 	src_data_18;
output 	src_payload70;
input 	readdata_82;
input 	d_writedata_22;
output 	src_payload71;
input 	readdata_222;
output 	src_payload72;
input 	readdata_72;
output 	src_payload73;
input 	readdata_62;
input 	readdata_201;
input 	d_writedata_20;
output 	src_payload74;
input 	readdata_191;
input 	d_writedata_19;
output 	src_payload75;
input 	readdata_04;
input 	read_0;
input 	av_readdata_0;
input 	readdata_05;
input 	counter_reg_bit_3;
input 	counter_reg_bit_0;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	b_full1;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	b_non_empty;
input 	counter_reg_bit_31;
input 	counter_reg_bit_21;
input 	counter_reg_bit_01;
input 	counter_reg_bit_11;
input 	counter_reg_bit_41;
input 	counter_reg_bit_51;
output 	src_payload76;
input 	readdata_113;
input 	av_readdata_1;
input 	readdata_114;
input 	readdata_210;
input 	av_readdata_2;
input 	readdata_213;
input 	readdata_33;
input 	av_readdata_3;
input 	readdata_34;
input 	readdata_43;
input 	av_readdata_4;
input 	readdata_44;
input 	readdata_53;
input 	av_readdata_5;
input 	readdata_54;
input 	readdata_63;
input 	av_readdata_6;
input 	readdata_64;
input 	readdata_73;
input 	av_readdata_7;
input 	readdata_74;
input 	readdata_83;
input 	readdata_92;
input 	readdata_102;
input 	ac;
input 	readdata_115;
input 	readdata_123;
input 	readdata_132;
input 	readdata_142;
input 	woverflow;
input 	readdata_152;
input 	rvalid;
input 	readdata_163;
input 	readdata_173;
output 	src_payload77;
output 	src_payload78;
output 	src_data_385;
output 	src_data_395;
output 	src_data_401;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_322;
output 	out_data_buffer_313;
output 	out_data_buffer_314;
output 	out_data_buffer_302;
output 	out_data_buffer_303;
output 	out_data_buffer_292;
output 	out_data_buffer_293;
output 	src_payload79;
output 	src_payload80;
output 	src_payload81;
input 	za_valid;
output 	out_data_buffer_02;
output 	out_data_buffer_110;
output 	src_payload82;
output 	out_data_buffer_210;
output 	src_payload83;
output 	src_payload84;
output 	src_payload85;
output 	src_data_331;
output 	src_payload86;
output 	src_payload87;
output 	src_data_341;
output 	src_payload88;
output 	src_payload89;
output 	src_payload90;
output 	src_payload91;
output 	src_payload92;
output 	src_payload93;
output 	src_payload94;
output 	src_payload95;
output 	src_data_351;
output 	src_payload96;
output 	src_payload97;
output 	src_payload98;
output 	src_payload99;
output 	src_payload100;
output 	src_payload101;
output 	src_payload102;
output 	src_payload103;
output 	src_payload104;
output 	src_payload105;
output 	src_payload106;
output 	src_payload107;
output 	src_payload108;
output 	src_payload109;
output 	src_payload110;
output 	src_payload111;
input 	za_data_0;
input 	za_data_1;
input 	za_data_2;
input 	za_data_3;
input 	za_data_4;
output 	src_payload112;
input 	za_data_11;
input 	za_data_13;
input 	za_data_16;
input 	za_data_12;
input 	za_data_5;
input 	za_data_14;
input 	za_data_15;
input 	za_data_21;
input 	za_data_18;
input 	za_data_17;
input 	za_data_31;
input 	za_data_30;
input 	za_data_29;
input 	za_data_28;
input 	za_data_27;
input 	za_data_26;
input 	za_data_25;
input 	za_data_10;
input 	za_data_24;
input 	za_data_9;
input 	za_data_23;
input 	za_data_8;
input 	za_data_22;
input 	za_data_7;
input 	za_data_6;
input 	za_data_20;
input 	za_data_19;
output 	src_payload113;
output 	src_payload114;
output 	src_payload115;
output 	src_payload116;
output 	src_payload117;
output 	src_payload118;
output 	src_payload119;
output 	src_payload120;
output 	src_payload121;
output 	src_payload122;
output 	src_payload123;
output 	src_payload124;
output 	src_payload125;
output 	src_payload126;
output 	src_payload127;
output 	src_payload128;
output 	src_payload129;
output 	src_payload130;
output 	src_payload131;
output 	src_payload132;
output 	src_payload133;
output 	src_payload134;
output 	src_payload135;
output 	src_payload136;
output 	src_payload137;
output 	src_payload138;
input 	av_ld_getting_data;
output 	m0_write;
output 	src_data_510;
output 	src_data_71;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \router|Equal8~4_combout ;
wire \router|Equal3~0_combout ;
wire \router|Equal0~0_combout ;
wire \router_001|Equal5~4_combout ;
wire \router_001|Equal0~0_combout ;
wire \router_001|Equal0~1_combout ;
wire \nios2_qsys_0_instruction_master_translator|read_accepted~q ;
wire \nios2_qsys_0_instruction_master_translator|uav_read~combout ;
wire \crosser_004|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_004|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \nios2_qsys_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][86]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \router|always1~0_combout ;
wire \router|src_channel[6]~5_combout ;
wire \router|src_channel[6]~6_combout ;
wire \router|Equal8~5_combout ;
wire \router|Equal2~3_combout ;
wire \router|src_channel[6]~7_combout ;
wire \router|Equal0~3_combout ;
wire \router|src_channel[9]~8_combout ;
wire \crosser_001|clock_xer|in_ready~0_combout ;
wire \cmd_demux|WideOr0~2_combout ;
wire \jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~2_combout ;
wire \router|Equal3~1_combout ;
wire \crosser|clock_xer|take_in_data~0_combout ;
wire \cmd_mux_004|saved_grant[0]~q ;
wire \router|Equal1~0_combout ;
wire \cmd_mux_005|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~9_combout ;
wire \cmd_mux_003|saved_grant[0]~q ;
wire \sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \router_001|Equal1~1_combout ;
wire \cmd_mux_003|saved_grant[1]~q ;
wire \cmd_mux_003|WideOr1~combout ;
wire \sysid_qsys_0_control_slave_agent|m0_write~0_combout ;
wire \sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~0_combout ;
wire \sysid_qsys_0_control_slave_agent|cp_ready~0_combout ;
wire \cmd_demux|WideOr0~10_combout ;
wire \rsp_mux_001|WideOr1~combout ;
wire \crosser_005|clock_xer|out_data_buffer[67]~q ;
wire \crosser_007|clock_xer|out_data_buffer[67]~q ;
wire \router_001|always1~1_combout ;
wire \cmd_mux_003|src_valid~0_combout ;
wire \router_001|Equal0~3_combout ;
wire \router_001|src_channel[6]~2_combout ;
wire \cmd_mux_009|saved_grant[1]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ;
wire \router_001|Equal6~0_combout ;
wire \router_001|Equal2~1_combout ;
wire \crosser_002|clock_xer|take_in_data~2_combout ;
wire \cmd_mux_005|saved_grant[1]~q ;
wire \router_001|Equal5~5_combout ;
wire \cmd_mux_004|saved_grant[1]~q ;
wire \router_001|src_channel[5]~3_combout ;
wire \crosser_003|clock_xer|in_ready~0_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \crosser_002|clock_xer|out_data_buffer[38]~q ;
wire \crosser|clock_xer|out_data_buffer[38]~q ;
wire \crosser_002|clock_xer|out_data_buffer[39]~q ;
wire \crosser|clock_xer|out_data_buffer[39]~q ;
wire \crosser_002|clock_xer|out_valid~combout ;
wire \crosser|clock_xer|out_data_toggle_flopped~q ;
wire \crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser|clock_xer|out_valid~combout ;
wire \crosser|clock_xer|out_data_buffer[67]~q ;
wire \ledg_s1_translator|wait_latency_counter[0]~0_combout ;
wire \ledr_s1_translator|wait_latency_counter[0]~0_combout ;
wire \sdram_s1_agent_rsp_fifo|mem_used[7]~q ;
wire \cmd_mux_006|saved_grant[0]~q ;
wire \crosser_003|clock_xer|out_valid~combout ;
wire \crosser_001|clock_xer|out_data_toggle_flopped~q ;
wire \crosser_001|clock_xer|in_to_out_synchronizer|dreg[0]~q ;
wire \crosser_001|clock_xer|out_valid~combout ;
wire \crosser_001|clock_xer|out_data_buffer[67]~q ;
wire \crosser_003|clock_xer|out_data_buffer[68]~q ;
wire \crosser_001|clock_xer|out_data_buffer[68]~q ;
wire \crosser_003|clock_xer|out_data_buffer[48]~q ;
wire \crosser_001|clock_xer|out_data_buffer[48]~q ;
wire \crosser_003|clock_xer|out_data_buffer[62]~q ;
wire \crosser_001|clock_xer|out_data_buffer[62]~q ;
wire \crosser_003|clock_xer|out_data_buffer[49]~q ;
wire \crosser_001|clock_xer|out_data_buffer[49]~q ;
wire \crosser_003|clock_xer|out_data_buffer[51]~q ;
wire \crosser_001|clock_xer|out_data_buffer[51]~q ;
wire \crosser_003|clock_xer|out_data_buffer[50]~q ;
wire \crosser_001|clock_xer|out_data_buffer[50]~q ;
wire \crosser_003|clock_xer|out_data_buffer[53]~q ;
wire \crosser_001|clock_xer|out_data_buffer[53]~q ;
wire \crosser_003|clock_xer|out_data_buffer[52]~q ;
wire \crosser_001|clock_xer|out_data_buffer[52]~q ;
wire \crosser_003|clock_xer|out_data_buffer[55]~q ;
wire \crosser_001|clock_xer|out_data_buffer[55]~q ;
wire \crosser_003|clock_xer|out_data_buffer[54]~q ;
wire \crosser_001|clock_xer|out_data_buffer[54]~q ;
wire \crosser_003|clock_xer|out_data_buffer[57]~q ;
wire \crosser_001|clock_xer|out_data_buffer[57]~q ;
wire \crosser_003|clock_xer|out_data_buffer[56]~q ;
wire \crosser_001|clock_xer|out_data_buffer[56]~q ;
wire \crosser_003|clock_xer|out_data_buffer[59]~q ;
wire \crosser_001|clock_xer|out_data_buffer[59]~q ;
wire \crosser_003|clock_xer|out_data_buffer[58]~q ;
wire \crosser_001|clock_xer|out_data_buffer[58]~q ;
wire \crosser_003|clock_xer|out_data_buffer[61]~q ;
wire \crosser_001|clock_xer|out_data_buffer[61]~q ;
wire \crosser_003|clock_xer|out_data_buffer[60]~q ;
wire \crosser_001|clock_xer|out_data_buffer[60]~q ;
wire \crosser_003|clock_xer|out_data_buffer[38]~q ;
wire \crosser_001|clock_xer|out_data_buffer[38]~q ;
wire \crosser_003|clock_xer|out_data_buffer[39]~q ;
wire \crosser_001|clock_xer|out_data_buffer[39]~q ;
wire \crosser_003|clock_xer|out_data_buffer[40]~q ;
wire \crosser_001|clock_xer|out_data_buffer[40]~q ;
wire \crosser_003|clock_xer|out_data_buffer[41]~q ;
wire \crosser_001|clock_xer|out_data_buffer[41]~q ;
wire \crosser_003|clock_xer|out_data_buffer[42]~q ;
wire \crosser_001|clock_xer|out_data_buffer[42]~q ;
wire \crosser_003|clock_xer|out_data_buffer[43]~q ;
wire \crosser_001|clock_xer|out_data_buffer[43]~q ;
wire \crosser_003|clock_xer|out_data_buffer[44]~q ;
wire \crosser_001|clock_xer|out_data_buffer[44]~q ;
wire \crosser_003|clock_xer|out_data_buffer[45]~q ;
wire \crosser_001|clock_xer|out_data_buffer[45]~q ;
wire \crosser_003|clock_xer|out_data_buffer[46]~q ;
wire \crosser_001|clock_xer|out_data_buffer[46]~q ;
wire \crosser_003|clock_xer|out_data_buffer[47]~q ;
wire \crosser_001|clock_xer|out_data_buffer[47]~q ;
wire \ledg_s1_translator|read_latency_shift_reg~0_combout ;
wire \ledr_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_mux_003|src_data[68]~combout ;
wire \sysid_qsys_0_control_slave_translator|read_latency_shift_reg~0_combout ;
wire \cmd_demux_001|src3_valid~0_combout ;
wire \nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ;
wire \sdram_pll_pll_slave_translator|read_latency_shift_reg~0_combout ;
wire \cmd_demux_001|src6_valid~0_combout ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem~1_combout ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \router|always1~2_combout ;
wire \cmd_mux_003|src_payload~0_combout ;
wire \crosser|clock_xer|out_data_buffer[31]~q ;
wire \audio_avalon_audio_slave_translator|waitrequest_reset_override~q ;
wire \crosser_002|clock_xer|out_data_buffer[107]~q ;
wire \crosser|clock_xer|out_data_buffer[107]~q ;
wire \cmd_mux|src_payload[0]~combout ;
wire \audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~0_combout ;
wire \audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~q ;
wire \audio_avalon_audio_slave_agent_rsp_fifo|mem[0][107]~q ;
wire \audio_avalon_audio_slave_translator|read_latency_shift_reg[0]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|mem_used[0]~q ;
wire \audio_avalon_audio_slave_agent|rp_valid~0_combout ;
wire \audio_avalon_audio_slave_agent_rsp_fifo|mem[0][86]~q ;
wire \audio_avalon_audio_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \crosser_005|clock_xer|in_data_toggle~q ;
wire \crosser_005|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_004|clock_xer|in_data_toggle~q ;
wire \crosser_004|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_005|clock_xer|take_in_data~0_combout ;
wire \rsp_demux|WideOr0~1_combout ;
wire \audio_avalon_audio_slave_agent|uncompressor|sink_ready~0_combout ;
wire \crosser|clock_xer|out_data_buffer[66]~q ;
wire \audio_avalon_audio_slave_agent|nonposted_write_endofpacket~1_combout ;
wire \crosser_002|clock_xer|out_data_buffer[68]~q ;
wire \crosser|clock_xer|out_data_buffer[68]~q ;
wire \crosser_003|clock_xer|out_data_buffer[107]~q ;
wire \crosser_001|clock_xer|out_data_buffer[107]~q ;
wire \cmd_mux_006|src_payload[0]~combout ;
wire \crosser_001|clock_xer|out_data_buffer[66]~q ;
wire \sdram_s1_agent|nonposted_write_endofpacket~0_combout ;
wire \sdram_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][107]~q ;
wire \sdram_s1_agent_rdata_fifo|out_valid~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][86]~q ;
wire \sdram_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \crosser_007|clock_xer|in_data_toggle~q ;
wire \crosser_007|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \crosser_006|clock_xer|in_data_toggle~q ;
wire \crosser_006|clock_xer|out_to_in_synchronizer|dreg[0]~q ;
wire \router_008|always0~0_combout ;
wire \rsp_demux_006|WideOr0~1_combout ;
wire \audio_avalon_audio_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \audio_avalon_audio_slave_agent|rp_valid~combout ;
wire \sdram_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \crosser_006|clock_xer|take_in_data~0_combout ;
wire \ledr_s1_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \crosser_006|clock_xer|out_data_buffer[0]~q ;
wire \crosser_004|clock_xer|out_data_buffer[0]~q ;
wire \ledg_s1_translator|av_readdata_pre[0]~q ;
wire \cmd_mux_003|src_data[38]~combout ;
wire \crosser|clock_xer|out_data_buffer[30]~q ;
wire \crosser_002|clock_xer|out_data_buffer[86]~q ;
wire \ledr_s1_translator|av_readdata_pre[1]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \crosser_006|clock_xer|out_data_buffer[1]~q ;
wire \ledg_s1_translator|av_readdata_pre[1]~q ;
wire \crosser_004|clock_xer|out_data_buffer[1]~q ;
wire \ledr_s1_translator|av_readdata_pre[2]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \crosser_006|clock_xer|out_data_buffer[2]~q ;
wire \ledg_s1_translator|av_readdata_pre[2]~q ;
wire \crosser_004|clock_xer|out_data_buffer[2]~q ;
wire \ledr_s1_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \crosser_006|clock_xer|out_data_buffer[3]~q ;
wire \ledg_s1_translator|av_readdata_pre[3]~q ;
wire \crosser_004|clock_xer|out_data_buffer[3]~q ;
wire \ledr_s1_translator|av_readdata_pre[4]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \crosser_006|clock_xer|out_data_buffer[4]~q ;
wire \ledg_s1_translator|av_readdata_pre[4]~q ;
wire \crosser_004|clock_xer|out_data_buffer[4]~q ;
wire \ledr_s1_translator|av_readdata_pre[5]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \crosser_006|clock_xer|out_data_buffer[5]~q ;
wire \ledg_s1_translator|av_readdata_pre[5]~q ;
wire \crosser_004|clock_xer|out_data_buffer[5]~q ;
wire \ledr_s1_translator|av_readdata_pre[6]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \crosser_006|clock_xer|out_data_buffer[6]~q ;
wire \ledg_s1_translator|av_readdata_pre[6]~q ;
wire \crosser_004|clock_xer|out_data_buffer[6]~q ;
wire \ledr_s1_translator|av_readdata_pre[7]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \crosser_006|clock_xer|out_data_buffer[7]~q ;
wire \ledg_s1_translator|av_readdata_pre[7]~q ;
wire \crosser_004|clock_xer|out_data_buffer[7]~q ;
wire \crosser_004|clock_xer|out_data_buffer[8]~q ;
wire \ledr_s1_translator|av_readdata_pre[8]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \crosser_006|clock_xer|out_data_buffer[8]~q ;
wire \ledr_s1_translator|av_readdata_pre[9]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \crosser_006|clock_xer|out_data_buffer[9]~q ;
wire \crosser_004|clock_xer|out_data_buffer[9]~q ;
wire \crosser_004|clock_xer|out_data_buffer[10]~q ;
wire \ledr_s1_translator|av_readdata_pre[10]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \crosser_006|clock_xer|out_data_buffer[10]~q ;
wire \crosser_006|clock_xer|out_data_buffer[11]~q ;
wire \crosser_004|clock_xer|out_data_buffer[11]~q ;
wire \ledr_s1_translator|av_readdata_pre[11]~q ;
wire \ledr_s1_translator|av_readdata_pre[12]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \crosser_006|clock_xer|out_data_buffer[12]~q ;
wire \crosser_004|clock_xer|out_data_buffer[12]~q ;
wire \ledr_s1_translator|av_readdata_pre[13]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \crosser_006|clock_xer|out_data_buffer[13]~q ;
wire \crosser_004|clock_xer|out_data_buffer[13]~q ;
wire \crosser_004|clock_xer|out_data_buffer[14]~q ;
wire \ledr_s1_translator|av_readdata_pre[14]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \crosser_006|clock_xer|out_data_buffer[14]~q ;
wire \ledr_s1_translator|av_readdata_pre[15]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \crosser_006|clock_xer|out_data_buffer[15]~q ;
wire \crosser_004|clock_xer|out_data_buffer[15]~q ;
wire \crosser_004|clock_xer|out_data_buffer[16]~q ;
wire \ledr_s1_translator|av_readdata_pre[16]~q ;
wire \crosser_006|clock_xer|out_data_buffer[16]~q ;
wire \crosser_004|clock_xer|out_data_buffer[17]~q ;
wire \crosser_006|clock_xer|out_data_buffer[17]~q ;
wire \ledr_s1_translator|av_readdata_pre[17]~q ;
wire \crosser_003|clock_xer|out_data_buffer[86]~q ;
wire \cmd_demux|WideOr0~11_combout ;
wire \crosser_001|clock_xer|out_data_buffer[0]~q ;
wire \crosser_001|clock_xer|out_data_buffer[1]~q ;
wire \crosser_001|clock_xer|out_data_buffer[2]~q ;
wire \crosser_001|clock_xer|out_data_buffer[3]~q ;
wire \crosser_001|clock_xer|out_data_buffer[4]~q ;
wire \crosser_001|clock_xer|out_data_buffer[5]~q ;
wire \crosser_001|clock_xer|out_data_buffer[6]~q ;
wire \crosser_001|clock_xer|out_data_buffer[7]~q ;
wire \crosser_001|clock_xer|out_data_buffer[8]~q ;
wire \crosser_001|clock_xer|out_data_buffer[9]~q ;
wire \crosser_001|clock_xer|out_data_buffer[10]~q ;
wire \crosser_001|clock_xer|out_data_buffer[11]~q ;
wire \crosser_001|clock_xer|out_data_buffer[12]~q ;
wire \crosser_001|clock_xer|out_data_buffer[13]~q ;
wire \crosser_001|clock_xer|out_data_buffer[14]~q ;
wire \crosser_001|clock_xer|out_data_buffer[15]~q ;
wire \crosser_001|clock_xer|out_data_buffer[16]~q ;
wire \crosser_001|clock_xer|out_data_buffer[17]~q ;
wire \crosser_001|clock_xer|out_data_buffer[18]~q ;
wire \crosser_001|clock_xer|out_data_buffer[19]~q ;
wire \crosser_001|clock_xer|out_data_buffer[20]~q ;
wire \crosser_001|clock_xer|out_data_buffer[21]~q ;
wire \crosser_001|clock_xer|out_data_buffer[22]~q ;
wire \crosser_001|clock_xer|out_data_buffer[23]~q ;
wire \crosser_001|clock_xer|out_data_buffer[24]~q ;
wire \crosser_001|clock_xer|out_data_buffer[25]~q ;
wire \crosser_001|clock_xer|out_data_buffer[26]~q ;
wire \crosser_001|clock_xer|out_data_buffer[27]~q ;
wire \crosser_001|clock_xer|out_data_buffer[28]~q ;
wire \crosser_001|clock_xer|out_data_buffer[29]~q ;
wire \crosser_001|clock_xer|out_data_buffer[30]~q ;
wire \crosser_001|clock_xer|out_data_buffer[31]~q ;
wire \crosser_004|clock_xer|out_data_buffer[23]~q ;
wire \crosser_006|clock_xer|out_data_buffer[23]~q ;
wire \crosser_004|clock_xer|out_data_buffer[22]~q ;
wire \crosser_006|clock_xer|out_data_buffer[22]~q ;
wire \crosser_006|clock_xer|out_data_buffer[21]~q ;
wire \crosser_004|clock_xer|out_data_buffer[21]~q ;
wire \crosser_006|clock_xer|out_data_buffer[20]~q ;
wire \crosser_004|clock_xer|out_data_buffer[20]~q ;
wire \crosser_006|clock_xer|out_data_buffer[19]~q ;
wire \crosser_004|clock_xer|out_data_buffer[19]~q ;
wire \crosser_004|clock_xer|out_data_buffer[18]~q ;
wire \crosser_006|clock_xer|out_data_buffer[18]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[0]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[0]~0_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[1]~1_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[1]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[2]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[2]~2_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[3]~3_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[3]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[4]~4_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[4]~q ;
wire \crosser|clock_xer|out_data_buffer[29]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[11]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[11]~5_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[13]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[13]~6_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[16]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[16]~7_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[12]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[12]~8_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[5]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[5]~9_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[14]~10_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[14]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[15]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[15]~11_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[21]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[21]~12_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[18]~13_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[18]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[17]~14_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[17]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[31]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[31]~15_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[30]~16_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[30]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[29]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[29]~17_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[28]~18_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[28]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[27]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[27]~19_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[26]~20_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[26]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[25]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[25]~21_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[10]~22_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[10]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[24]~23_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[24]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[9]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[9]~24_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[23]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[23]~25_combout ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[8]~26_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[8]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[22]~27_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[22]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[7]~28_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[7]~q ;
wire \sdram_s1_agent_rdata_fifo|out_payload[6]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[6]~29_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[20]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[20]~30_combout ;
wire \sdram_s1_agent_rdata_fifo|out_payload[19]~q ;
wire \audio_avalon_audio_slave_agent_rdata_fifo|out_data[19]~31_combout ;
wire \crosser|clock_xer|out_data_buffer[28]~q ;
wire \crosser|clock_xer|out_data_buffer[27]~q ;
wire \crosser|clock_xer|out_data_buffer[26]~q ;
wire \crosser|clock_xer|out_data_buffer[25]~q ;
wire \crosser|clock_xer|out_data_buffer[24]~q ;
wire \crosser|clock_xer|out_data_buffer[23]~q ;
wire \crosser|clock_xer|out_data_buffer[22]~q ;
wire \crosser|clock_xer|out_data_buffer[21]~q ;
wire \crosser|clock_xer|out_data_buffer[20]~q ;
wire \crosser|clock_xer|out_data_buffer[19]~q ;
wire \crosser|clock_xer|out_data_buffer[18]~q ;
wire \crosser|clock_xer|out_data_buffer[17]~q ;
wire \crosser|clock_xer|out_data_buffer[16]~q ;
wire \crosser|clock_xer|out_data_buffer[15]~q ;
wire \crosser|clock_xer|out_data_buffer[14]~q ;
wire \crosser|clock_xer|out_data_buffer[13]~q ;
wire \crosser|clock_xer|out_data_buffer[12]~q ;
wire \crosser|clock_xer|out_data_buffer[11]~q ;
wire \crosser|clock_xer|out_data_buffer[10]~q ;
wire \crosser|clock_xer|out_data_buffer[9]~q ;
wire \crosser|clock_xer|out_data_buffer[8]~q ;
wire \crosser|clock_xer|out_data_buffer[7]~q ;
wire \crosser|clock_xer|out_data_buffer[6]~q ;
wire \crosser|clock_xer|out_data_buffer[5]~q ;
wire \crosser|clock_xer|out_data_buffer[4]~q ;
wire \cmd_demux_001|src4_valid~2_combout ;


final_project_soc_altera_avalon_sc_fifo_9 sdram_s1_agent_rdata_fifo(
	.clk(wire_pll7_clk_0),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\sdram_s1_agent_rsp_fifo|mem[0][107]~q ),
	.out_valid1(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.WideOr0(\rsp_demux_006|WideOr0~1_combout ),
	.out_payload_0(\sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.out_payload_1(\sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.out_payload_2(\sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.out_payload_3(\sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.out_payload_4(\sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.out_payload_11(\sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.out_payload_13(\sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.out_payload_16(\sdram_s1_agent_rdata_fifo|out_payload[16]~q ),
	.out_payload_12(\sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.out_payload_5(\sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.out_payload_14(\sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.out_payload_15(\sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.out_payload_21(\sdram_s1_agent_rdata_fifo|out_payload[21]~q ),
	.out_payload_18(\sdram_s1_agent_rdata_fifo|out_payload[18]~q ),
	.out_payload_17(\sdram_s1_agent_rdata_fifo|out_payload[17]~q ),
	.out_payload_31(\sdram_s1_agent_rdata_fifo|out_payload[31]~q ),
	.out_payload_30(\sdram_s1_agent_rdata_fifo|out_payload[30]~q ),
	.out_payload_29(\sdram_s1_agent_rdata_fifo|out_payload[29]~q ),
	.out_payload_28(\sdram_s1_agent_rdata_fifo|out_payload[28]~q ),
	.out_payload_27(\sdram_s1_agent_rdata_fifo|out_payload[27]~q ),
	.out_payload_26(\sdram_s1_agent_rdata_fifo|out_payload[26]~q ),
	.out_payload_25(\sdram_s1_agent_rdata_fifo|out_payload[25]~q ),
	.out_payload_10(\sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.out_payload_24(\sdram_s1_agent_rdata_fifo|out_payload[24]~q ),
	.out_payload_9(\sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.out_payload_23(\sdram_s1_agent_rdata_fifo|out_payload[23]~q ),
	.out_payload_8(\sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.out_payload_22(\sdram_s1_agent_rdata_fifo|out_payload[22]~q ),
	.out_payload_7(\sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.out_payload_6(\sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.out_payload_20(\sdram_s1_agent_rdata_fifo|out_payload[20]~q ),
	.out_payload_19(\sdram_s1_agent_rdata_fifo|out_payload[19]~q ),
	.za_valid(za_valid),
	.za_data_0(za_data_0),
	.za_data_1(za_data_1),
	.za_data_2(za_data_2),
	.za_data_3(za_data_3),
	.za_data_4(za_data_4),
	.za_data_11(za_data_11),
	.za_data_13(za_data_13),
	.za_data_16(za_data_16),
	.za_data_12(za_data_12),
	.za_data_5(za_data_5),
	.za_data_14(za_data_14),
	.za_data_15(za_data_15),
	.za_data_21(za_data_21),
	.za_data_18(za_data_18),
	.za_data_17(za_data_17),
	.za_data_31(za_data_31),
	.za_data_30(za_data_30),
	.za_data_29(za_data_29),
	.za_data_28(za_data_28),
	.za_data_27(za_data_27),
	.za_data_26(za_data_26),
	.za_data_25(za_data_25),
	.za_data_10(za_data_10),
	.za_data_24(za_data_24),
	.za_data_9(za_data_9),
	.za_data_23(za_data_23),
	.za_data_8(za_data_8),
	.za_data_22(za_data_22),
	.za_data_7(za_data_7),
	.za_data_6(za_data_6),
	.za_data_20(za_data_20),
	.za_data_19(za_data_19));

final_project_soc_altera_avalon_sc_fifo_10 sdram_s1_agent_rsp_fifo(
	.clk(wire_pll7_clk_0),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.last_cycle(last_cycle1),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.saved_grant_1(saved_grant_11),
	.WideOr1(WideOr14),
	.out_data_buffer_67(\crosser_001|clock_xer|out_data_buffer[67]~q ),
	.src_data_68(src_data_681),
	.nonposted_write_endofpacket(\sdram_s1_agent|nonposted_write_endofpacket~0_combout ),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\sdram_s1_agent_rsp_fifo|mem[0][107]~q ),
	.out_valid(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.WideOr0(\rsp_demux_006|WideOr0~1_combout ),
	.mem_67_0(\sdram_s1_agent_rsp_fifo|mem[0][67]~q ),
	.out_data_buffer_86(\crosser_003|clock_xer|out_data_buffer[86]~q ));

final_project_soc_altera_merlin_slave_agent_8 sdram_s1_agent(
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.WideOr1(WideOr14),
	.out_data_buffer_67(\crosser_001|clock_xer|out_data_buffer[67]~q ),
	.src_payload(src_payload3),
	.src_payload_0(\cmd_mux_006|src_payload[0]~combout ),
	.out_data_buffer_66(\crosser_001|clock_xer|out_data_buffer[66]~q ),
	.nonposted_write_endofpacket(\sdram_s1_agent|nonposted_write_endofpacket~0_combout ),
	.m0_write(m0_write));

final_project_soc_altera_avalon_sc_fifo_8 sdram_pll_pll_slave_agent_rsp_fifo(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.uav_read1(uav_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.mem_86_0(mem_86_01),
	.mem_68_0(mem_68_01),
	.mem_67_0(mem_67_03),
	.rst1(rst1),
	.saved_grant_0(\cmd_mux_005|saved_grant[0]~q ),
	.mem_used_1(mem_used_15),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.WideOr1(WideOr13),
	.mem(mem),
	.mem1(mem1),
	.read_latency_shift_reg(\sdram_pll_pll_slave_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_avalon_sc_fifo_6 nios2_qsys_0_debug_mem_slave_agent_rsp_fifo(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.uav_read1(uav_read),
	.read_latency_shift_reg_0(\nios2_qsys_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(mem_67_02),
	.saved_grant_0(\cmd_mux_004|saved_grant[0]~q ),
	.waitrequest(waitrequest1),
	.mem_used_1(mem_used_14),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.mem(\nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.local_read(local_read),
	.mem1(mem2),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_agent_5 nios2_qsys_0_debug_mem_slave_agent(
	.WideOr1(WideOr15),
	.mem(\nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.local_read(local_read));

final_project_soc_altera_avalon_sc_fifo_11 sysid_qsys_0_control_slave_agent_rsp_fifo(
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(mem_67_01),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.WideOr1(\cmd_mux_003|WideOr1~combout ),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ),
	.src_data_68(\cmd_mux_003|src_data[68]~combout ),
	.read_latency_shift_reg(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_agent_9 sysid_qsys_0_control_slave_agent(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.rst1(rst1),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\sysid_qsys_0_control_slave_agent|m0_write~0_combout ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~0_combout ),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ));

final_project_soc_altera_avalon_sc_fifo_3 jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo(
	.d_read(d_read),
	.d_write(d_write),
	.read_accepted(read_accepted),
	.write_accepted(write_accepted),
	.reset(r_sync_rst),
	.uav_read(uav_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_67_0(mem_67_04),
	.Equal2(\router|Equal2~3_combout ),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~2_combout ),
	.clk(clk_clk));

final_project_soc_altera_avalon_sc_fifo_2 audio_config_avalon_av_config_slave_agent_rsp_fifo(
	.saved_grant_1(saved_grant_1),
	.saved_grant_0(saved_grant_0),
	.uav_write(uav_write),
	.mem_used_1(mem_used_1),
	.reset(r_sync_rst),
	.WideOr1(WideOr1),
	.src_data_68(src_data_68),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.waitrequest(waitrequest2),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_agent_1 audio_config_avalon_av_config_slave_agent(
	.mem_used_1(mem_used_1),
	.WideOr1(WideOr1),
	.src_data_68(src_data_68),
	.m0_read1(m0_read));

final_project_soc_altera_avalon_sc_fifo audio_avalon_audio_slave_agent_rdata_fifo(
	.clk(clk_0),
	.readdata_0(readdata_02),
	.readdata_1(readdata_12),
	.readdata_2(readdata_22),
	.readdata_3(readdata_31),
	.readdata_4(readdata_4),
	.readdata_11(readdata_111),
	.readdata_13(readdata_13),
	.readdata_16(readdata_161),
	.readdata_12(readdata_121),
	.readdata_5(readdata_5),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_21(readdata_211),
	.readdata_18(readdata_18),
	.readdata_17(readdata_171),
	.readdata_31(readdata_311),
	.readdata_30(readdata_30),
	.readdata_29(readdata_29),
	.readdata_28(readdata_28),
	.readdata_27(readdata_27),
	.readdata_26(readdata_26),
	.readdata_25(readdata_25),
	.readdata_10(readdata_10),
	.readdata_24(readdata_24),
	.readdata_9(readdata_9),
	.readdata_23(readdata_23),
	.readdata_8(readdata_81),
	.readdata_22(readdata_221),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.reset(altera_reset_synchronizer_int_chain_out),
	.mem_used_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][107]~q ),
	.read_latency_shift_reg_0(\audio_avalon_audio_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\audio_avalon_audio_slave_agent_rdata_fifo|mem_used[0]~q ),
	.rp_valid(\audio_avalon_audio_slave_agent|rp_valid~0_combout ),
	.WideOr0(\rsp_demux|WideOr0~1_combout ),
	.out_data_0(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_11(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[11]~5_combout ),
	.out_data_13(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[13]~6_combout ),
	.out_data_16(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[16]~7_combout ),
	.out_data_12(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[12]~8_combout ),
	.out_data_5(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[5]~9_combout ),
	.out_data_14(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[14]~10_combout ),
	.out_data_15(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[15]~11_combout ),
	.out_data_21(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[21]~12_combout ),
	.out_data_18(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[18]~13_combout ),
	.out_data_17(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[17]~14_combout ),
	.out_data_31(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[31]~15_combout ),
	.out_data_30(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[30]~16_combout ),
	.out_data_29(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[29]~17_combout ),
	.out_data_28(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[28]~18_combout ),
	.out_data_27(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[27]~19_combout ),
	.out_data_26(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[26]~20_combout ),
	.out_data_25(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[25]~21_combout ),
	.out_data_10(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[10]~22_combout ),
	.out_data_24(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[24]~23_combout ),
	.out_data_9(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[9]~24_combout ),
	.out_data_23(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[23]~25_combout ),
	.out_data_8(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[8]~26_combout ),
	.out_data_22(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[22]~27_combout ),
	.out_data_7(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[7]~28_combout ),
	.out_data_6(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[6]~29_combout ),
	.out_data_20(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[20]~30_combout ),
	.out_data_19(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[19]~31_combout ));

final_project_soc_altera_avalon_sc_fifo_1 audio_avalon_audio_slave_agent_rsp_fifo(
	.clk(clk_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.saved_grant_0(saved_grant_02),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.WideOr1(WideOr12),
	.mem_used_1(mem_used_17),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.waitrequest_reset_override(\audio_avalon_audio_slave_translator|waitrequest_reset_override~q ),
	.mem_used_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~0_combout ),
	.mem_used_01(\audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][107]~q ),
	.rp_valid(\audio_avalon_audio_slave_agent|rp_valid~0_combout ),
	.mem_86_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][68]~q ),
	.WideOr0(\rsp_demux|WideOr0~1_combout ),
	.sink_ready(\audio_avalon_audio_slave_agent|uncompressor|sink_ready~0_combout ),
	.nonposted_write_endofpacket(\audio_avalon_audio_slave_agent|nonposted_write_endofpacket~1_combout ),
	.src_data_68(src_data_682),
	.mem_67_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][67]~q ),
	.out_data_buffer_86(\crosser_002|clock_xer|out_data_buffer[86]~q ));

final_project_soc_altera_merlin_slave_agent audio_avalon_audio_slave_agent(
	.saved_grant_0(saved_grant_02),
	.WideOr1(WideOr12),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.nonposted_write_endofpacket(nonposted_write_endofpacket),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.mem_used_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][107]~q ),
	.read_latency_shift_reg_0(\audio_avalon_audio_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\audio_avalon_audio_slave_agent_rdata_fifo|mem_used[0]~q ),
	.rp_valid1(\audio_avalon_audio_slave_agent|rp_valid~0_combout ),
	.WideOr0(\rsp_demux|WideOr0~1_combout ),
	.rf_sink_ready(\audio_avalon_audio_slave_agent|uncompressor|sink_ready~0_combout ),
	.out_data_buffer_66(\crosser|clock_xer|out_data_buffer[66]~q ),
	.nonposted_write_endofpacket1(\audio_avalon_audio_slave_agent|nonposted_write_endofpacket~1_combout ),
	.rp_valid2(\audio_avalon_audio_slave_agent|rp_valid~combout ));

final_project_soc_altera_merlin_master_agent_1 nios2_qsys_0_instruction_master_agent(
	.mem_67_0(mem_67_0),
	.mem_67_01(mem_67_01),
	.mem_67_02(mem_67_02),
	.mem_67_03(mem_67_03),
	.mem_67_04(mem_67_06),
	.src1_valid(src1_valid1),
	.src1_valid1(src1_valid2),
	.src1_valid2(src1_valid3),
	.src_payload(src_payload1),
	.src_payload1(src_payload2),
	.out_valid(out_valid2),
	.out_valid1(out_valid3),
	.WideOr1(\rsp_mux_001|WideOr1~combout ),
	.out_data_buffer_67(\crosser_005|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_671(\crosser_007|clock_xer|out_data_buffer[67]~q ),
	.av_readdatavalid(av_readdatavalid));

final_project_soc_altera_merlin_master_agent nios2_qsys_0_data_master_agent(
	.d_read(d_read),
	.d_write(d_write),
	.read_accepted(read_accepted),
	.write_accepted(write_accepted),
	.cp_valid1(cp_valid));

final_project_soc_altera_merlin_slave_translator_6 onchip_memory2_0_s1_translator(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.rst1(rst1),
	.mem_used_1(mem_used_16),
	.WideOr1(WideOr16),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~1_combout ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_3 ledg_s1_translator(
	.cp_valid(cp_valid),
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.always0(always0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.uav_read(uav_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.rst1(rst1),
	.wait_latency_counter_01(\ledg_s1_translator|wait_latency_counter[0]~0_combout ),
	.read_latency_shift_reg(\ledg_s1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(\ledg_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\ledg_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\ledg_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\ledg_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\ledg_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\ledg_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\ledg_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\ledg_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_74,readdata_64,readdata_54,readdata_44,readdata_34,readdata_213,readdata_114,readdata_05}),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_4 ledr_s1_translator(
	.cp_valid(cp_valid),
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.always0(always01),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.uav_read(uav_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.rst1(rst1),
	.wait_latency_counter_01(\ledr_s1_translator|wait_latency_counter[0]~0_combout ),
	.read_latency_shift_reg(\ledr_s1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(\ledr_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\ledr_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\ledr_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\ledr_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\ledr_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\ledr_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\ledr_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\ledr_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\ledr_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\ledr_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\ledr_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\ledr_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\ledr_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\ledr_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\ledr_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\ledr_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\ledr_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\ledr_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_173,readdata_163,readdata_152,readdata_142,readdata_132,readdata_123,readdata_115,readdata_102,readdata_92,readdata_83,readdata_73,readdata_63,readdata_53,readdata_43,readdata_33,readdata_210,readdata_113,readdata_04}),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_7 sdram_pll_pll_slave_translator(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.rst1(rst1),
	.mem_used_1(mem_used_15),
	.WideOr1(WideOr13),
	.mem(mem1),
	.read_latency_shift_reg(\sdram_pll_pll_slave_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(av_readdata_pre_01),
	.av_readdata_pre_1(av_readdata_pre_11),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_110,readdata_03}),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_5 nios2_qsys_0_debug_mem_slave_translator(
	.av_readdata({readdata_312,readdata_301,readdata_291,readdata_281,readdata_271,readdata_261,readdata_251,readdata_241,readdata_231,readdata_222,readdata_212,readdata_201,readdata_191,readdata_181,readdata_172,readdata_162,readdata_151,readdata_141,readdata_131,readdata_122,readdata_112,
readdata_101,readdata_91,readdata_82,readdata_72,readdata_62,readdata_52,readdata_42,readdata_3,readdata_21,readdata_11,readdata_01}),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\nios2_qsys_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.rst1(rst1),
	.waitrequest(waitrequest1),
	.mem_used_1(mem_used_14),
	.local_read(local_read),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_11(av_readdata_pre_111),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_30(av_readdata_pre_301),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_19(av_readdata_pre_19),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_9 sysid_qsys_0_control_slave_translator(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.rst1(rst1),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr1(\cmd_mux_003|WideOr1~combout ),
	.m0_write(\sysid_qsys_0_control_slave_agent|m0_write~0_combout ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~0_combout ),
	.src_data_68(\cmd_mux_003|src_data[68]~combout ),
	.read_latency_shift_reg(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg~0_combout ),
	.src_payload(\cmd_mux_003|src_payload~0_combout ),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata({gnd,\cmd_mux_003|src_data[38]~combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_2 jtag_uart_0_avalon_jtag_slave_translator(
	.av_readdata_pre_16(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_22(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.reset(r_sync_rst),
	.Equal2(Equal2),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.rst1(rst1),
	.Equal21(Equal22),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~2_combout ),
	.av_readdata_pre_0(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,av_readdata_7,av_readdata_6,av_readdata_5,av_readdata_4,av_readdata_3,av_readdata_2,av_readdata_1,av_readdata_0}),
	.av_readdata_pre_1(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_12(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.b_full(b_full),
	.read_0(read_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full1(b_full1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_31(counter_reg_bit_31),
	.counter_reg_bit_21(counter_reg_bit_21),
	.counter_reg_bit_01(counter_reg_bit_01),
	.counter_reg_bit_11(counter_reg_bit_11),
	.counter_reg_bit_41(counter_reg_bit_41),
	.counter_reg_bit_51(counter_reg_bit_51),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator_1 audio_config_avalon_av_config_slave_translator(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.rst1(rst1),
	.waitrequest(waitrequest2),
	.m0_read(m0_read),
	.clk(clk_clk));

final_project_soc_altera_merlin_slave_translator audio_avalon_audio_slave_translator(
	.clk(clk_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr1(WideOr12),
	.mem_used_1(mem_used_17),
	.waitrequest_reset_override1(\audio_avalon_audio_slave_translator|waitrequest_reset_override~q ),
	.read_latency_shift_reg_0(\audio_avalon_audio_slave_translator|read_latency_shift_reg[0]~q ),
	.src_data_68(src_data_682));

final_project_soc_altera_merlin_master_translator_1 nios2_qsys_0_instruction_master_translator(
	.saved_grant_1(saved_grant_1),
	.F_pc_5(F_pc_5),
	.i_read(i_read),
	.read_accepted1(\nios2_qsys_0_instruction_master_translator|read_accepted~q ),
	.uav_read1(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.F_pc_2(F_pc_2),
	.mem_used_1(mem_used_1),
	.reset(r_sync_rst),
	.rst1(rst1),
	.waitrequest(waitrequest1),
	.mem_used_11(mem_used_14),
	.mem_used_12(mem_used_15),
	.waitrequest1(waitrequest2),
	.mem_used_13(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.Equal1(\router_001|Equal1~1_combout ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~0_combout ),
	.av_readdatavalid(av_readdatavalid),
	.src_valid(\cmd_mux_003|src_valid~0_combout ),
	.Equal0(\router_001|Equal0~3_combout ),
	.src_channel_6(\router_001|src_channel[6]~2_combout ),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ),
	.Equal6(\router_001|Equal6~0_combout ),
	.Equal2(\router_001|Equal2~1_combout ),
	.take_in_data(\crosser_002|clock_xer|take_in_data~2_combout ),
	.saved_grant_11(\cmd_mux_005|saved_grant[1]~q ),
	.Equal5(\router_001|Equal5~5_combout ),
	.saved_grant_12(\cmd_mux_004|saved_grant[1]~q ),
	.src_channel_5(\router_001|src_channel[5]~3_combout ),
	.in_ready(\crosser_003|clock_xer|in_ready~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_merlin_master_translator nios2_qsys_0_data_master_translator(
	.d_read(d_read),
	.d_write(d_write),
	.read_accepted1(read_accepted),
	.write_accepted1(write_accepted),
	.cp_valid(cp_valid),
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.uav_read(uav_read),
	.rst1(rst1),
	.WideOr0(\cmd_demux|WideOr0~9_combout ),
	.WideOr01(\cmd_demux|WideOr0~10_combout ),
	.av_waitrequest(nios2_qsys_0_data_master_waitrequest),
	.av_ld_getting_data(av_ld_getting_data),
	.clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001 rsp_demux_001(
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid1));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux rsp_demux(
	.mem_86_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][68]~q ),
	.in_data_toggle(\crosser_005|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_005|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.in_data_toggle1(\crosser_004|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_004|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.take_in_data(\crosser_005|clock_xer|take_in_data~0_combout ),
	.WideOr0(\rsp_demux|WideOr0~1_combout ));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_6 cmd_mux_009(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_31(d_writedata_31),
	.d_writedata_30(d_writedata_30),
	.d_writedata_29(d_writedata_29),
	.d_writedata_28(d_writedata_28),
	.d_writedata_27(d_writedata_27),
	.d_writedata_26(d_writedata_26),
	.d_writedata_25(d_writedata_25),
	.d_writedata_24(d_writedata_24),
	.cp_valid(cp_valid),
	.d_writedata_0(d_writedata_0),
	.d_byteenable_0(d_byteenable_0),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.Equal0(Equal0),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.rst1(rst1),
	.src_channel_6(\router|src_channel[6]~5_combout ),
	.src_channel_61(\router|src_channel[6]~6_combout ),
	.Equal8(\router|Equal8~5_combout ),
	.Equal2(\router|Equal2~3_combout ),
	.src_channel_9(\router|src_channel[9]~8_combout ),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_16),
	.saved_grant_1(\cmd_mux_009|saved_grant[1]~q ),
	.src6_valid(\cmd_demux_001|src6_valid~0_combout ),
	.WideOr11(WideOr16),
	.d_byteenable_2(d_byteenable_2),
	.src_payload(src_payload11),
	.src_data_38(src_data_384),
	.src_data_39(src_data_394),
	.src_data_32(src_data_321),
	.src_payload1(src_payload12),
	.src_payload2(src_payload13),
	.src_payload3(src_payload14),
	.src_payload4(src_payload15),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_3(d_byteenable_3),
	.src_payload5(src_payload49),
	.src_data_33(src_data_33),
	.src_payload6(src_payload50),
	.src_payload7(src_payload51),
	.src_data_34(src_data_34),
	.src_payload8(src_payload52),
	.src_payload9(src_payload53),
	.src_payload10(src_payload54),
	.src_payload11(src_payload55),
	.d_writedata_21(d_writedata_21),
	.src_payload12(src_payload56),
	.d_writedata_18(d_writedata_18),
	.src_payload13(src_payload57),
	.src_payload14(src_payload58),
	.src_payload15(src_payload59),
	.src_data_35(src_data_35),
	.src_payload16(src_payload60),
	.src_payload17(src_payload61),
	.src_payload18(src_payload62),
	.src_payload19(src_payload63),
	.src_payload20(src_payload64),
	.src_payload21(src_payload65),
	.src_payload22(src_payload66),
	.src_payload23(src_payload67),
	.src_payload24(src_payload68),
	.d_writedata_23(d_writedata_23),
	.src_payload25(src_payload69),
	.src_payload26(src_payload70),
	.d_writedata_22(d_writedata_22),
	.src_payload27(src_payload71),
	.src_payload28(src_payload72),
	.src_payload29(src_payload73),
	.d_writedata_20(d_writedata_20),
	.src_payload30(src_payload74),
	.d_writedata_19(d_writedata_19),
	.src_payload31(src_payload75),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_5 cmd_mux_006(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.mem_used_7(\sdram_s1_agent_rsp_fifo|mem_used[7]~q ),
	.last_cycle(last_cycle1),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.saved_grant_1(saved_grant_11),
	.out_valid(\crosser_003|clock_xer|out_valid~combout ),
	.out_data_toggle_flopped(\crosser_001|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_001|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid1(\crosser_001|clock_xer|out_valid~combout ),
	.WideOr11(WideOr14),
	.out_data_buffer_67(\crosser_001|clock_xer|out_data_buffer[67]~q ),
	.src_payload(src_payload3),
	.out_data_buffer_68(\crosser_003|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_681(\crosser_001|clock_xer|out_data_buffer[68]~q ),
	.src_data_68(src_data_681),
	.out_data_buffer_48(\crosser_003|clock_xer|out_data_buffer[48]~q ),
	.out_data_buffer_481(\crosser_001|clock_xer|out_data_buffer[48]~q ),
	.src_data_48(src_data_48),
	.out_data_buffer_62(\crosser_003|clock_xer|out_data_buffer[62]~q ),
	.out_data_buffer_621(\crosser_001|clock_xer|out_data_buffer[62]~q ),
	.src_data_62(src_data_62),
	.out_data_buffer_49(\crosser_003|clock_xer|out_data_buffer[49]~q ),
	.out_data_buffer_491(\crosser_001|clock_xer|out_data_buffer[49]~q ),
	.src_data_49(src_data_49),
	.out_data_buffer_51(\crosser_003|clock_xer|out_data_buffer[51]~q ),
	.out_data_buffer_511(\crosser_001|clock_xer|out_data_buffer[51]~q ),
	.src_data_51(src_data_51),
	.out_data_buffer_50(\crosser_003|clock_xer|out_data_buffer[50]~q ),
	.out_data_buffer_501(\crosser_001|clock_xer|out_data_buffer[50]~q ),
	.src_data_50(src_data_50),
	.out_data_buffer_53(\crosser_003|clock_xer|out_data_buffer[53]~q ),
	.out_data_buffer_531(\crosser_001|clock_xer|out_data_buffer[53]~q ),
	.src_data_53(src_data_53),
	.out_data_buffer_52(\crosser_003|clock_xer|out_data_buffer[52]~q ),
	.out_data_buffer_521(\crosser_001|clock_xer|out_data_buffer[52]~q ),
	.src_data_52(src_data_52),
	.out_data_buffer_55(\crosser_003|clock_xer|out_data_buffer[55]~q ),
	.out_data_buffer_551(\crosser_001|clock_xer|out_data_buffer[55]~q ),
	.src_data_55(src_data_55),
	.out_data_buffer_54(\crosser_003|clock_xer|out_data_buffer[54]~q ),
	.out_data_buffer_541(\crosser_001|clock_xer|out_data_buffer[54]~q ),
	.src_data_54(src_data_54),
	.out_data_buffer_57(\crosser_003|clock_xer|out_data_buffer[57]~q ),
	.out_data_buffer_571(\crosser_001|clock_xer|out_data_buffer[57]~q ),
	.src_data_57(src_data_57),
	.out_data_buffer_56(\crosser_003|clock_xer|out_data_buffer[56]~q ),
	.out_data_buffer_561(\crosser_001|clock_xer|out_data_buffer[56]~q ),
	.src_data_56(src_data_56),
	.out_data_buffer_59(\crosser_003|clock_xer|out_data_buffer[59]~q ),
	.out_data_buffer_591(\crosser_001|clock_xer|out_data_buffer[59]~q ),
	.src_data_59(src_data_59),
	.out_data_buffer_58(\crosser_003|clock_xer|out_data_buffer[58]~q ),
	.out_data_buffer_581(\crosser_001|clock_xer|out_data_buffer[58]~q ),
	.src_data_58(src_data_58),
	.out_data_buffer_61(\crosser_003|clock_xer|out_data_buffer[61]~q ),
	.out_data_buffer_611(\crosser_001|clock_xer|out_data_buffer[61]~q ),
	.src_data_61(src_data_61),
	.out_data_buffer_60(\crosser_003|clock_xer|out_data_buffer[60]~q ),
	.out_data_buffer_601(\crosser_001|clock_xer|out_data_buffer[60]~q ),
	.src_data_60(src_data_60),
	.out_data_buffer_38(\crosser_003|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_381(\crosser_001|clock_xer|out_data_buffer[38]~q ),
	.src_data_38(src_data_383),
	.out_data_buffer_39(\crosser_003|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_391(\crosser_001|clock_xer|out_data_buffer[39]~q ),
	.src_data_39(src_data_393),
	.out_data_buffer_40(\crosser_003|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_401(\crosser_001|clock_xer|out_data_buffer[40]~q ),
	.src_data_40(src_data_40),
	.out_data_buffer_41(\crosser_003|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_411(\crosser_001|clock_xer|out_data_buffer[41]~q ),
	.src_data_41(src_data_41),
	.out_data_buffer_42(\crosser_003|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_421(\crosser_001|clock_xer|out_data_buffer[42]~q ),
	.src_data_42(src_data_42),
	.out_data_buffer_43(\crosser_003|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_431(\crosser_001|clock_xer|out_data_buffer[43]~q ),
	.src_data_43(src_data_43),
	.out_data_buffer_44(\crosser_003|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_441(\crosser_001|clock_xer|out_data_buffer[44]~q ),
	.src_data_44(src_data_44),
	.out_data_buffer_45(\crosser_003|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_451(\crosser_001|clock_xer|out_data_buffer[45]~q ),
	.src_data_45(src_data_45),
	.out_data_buffer_46(\crosser_003|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_461(\crosser_001|clock_xer|out_data_buffer[46]~q ),
	.src_data_46(src_data_46),
	.out_data_buffer_47(\crosser_003|clock_xer|out_data_buffer[47]~q ),
	.out_data_buffer_471(\crosser_001|clock_xer|out_data_buffer[47]~q ),
	.src_data_47(src_data_47),
	.out_data_buffer_107(\crosser_003|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_1071(\crosser_001|clock_xer|out_data_buffer[107]~q ),
	.src_payload_0(\cmd_mux_006|src_payload[0]~combout ),
	.out_data_buffer_0(\crosser_001|clock_xer|out_data_buffer[0]~q ),
	.src_payload1(src_payload17),
	.out_data_buffer_1(\crosser_001|clock_xer|out_data_buffer[1]~q ),
	.src_payload2(src_payload18),
	.out_data_buffer_2(\crosser_001|clock_xer|out_data_buffer[2]~q ),
	.src_payload3(src_payload19),
	.out_data_buffer_3(\crosser_001|clock_xer|out_data_buffer[3]~q ),
	.src_payload4(src_payload20),
	.out_data_buffer_4(\crosser_001|clock_xer|out_data_buffer[4]~q ),
	.src_payload5(src_payload21),
	.out_data_buffer_5(\crosser_001|clock_xer|out_data_buffer[5]~q ),
	.src_payload6(src_payload22),
	.out_data_buffer_6(\crosser_001|clock_xer|out_data_buffer[6]~q ),
	.src_payload7(src_payload23),
	.out_data_buffer_7(\crosser_001|clock_xer|out_data_buffer[7]~q ),
	.src_payload8(src_payload24),
	.out_data_buffer_8(\crosser_001|clock_xer|out_data_buffer[8]~q ),
	.src_payload9(src_payload25),
	.out_data_buffer_9(\crosser_001|clock_xer|out_data_buffer[9]~q ),
	.src_payload10(src_payload26),
	.out_data_buffer_10(\crosser_001|clock_xer|out_data_buffer[10]~q ),
	.src_payload11(src_payload27),
	.out_data_buffer_11(\crosser_001|clock_xer|out_data_buffer[11]~q ),
	.src_payload12(src_payload28),
	.out_data_buffer_12(\crosser_001|clock_xer|out_data_buffer[12]~q ),
	.src_payload13(src_payload29),
	.out_data_buffer_13(\crosser_001|clock_xer|out_data_buffer[13]~q ),
	.src_payload14(src_payload30),
	.out_data_buffer_14(\crosser_001|clock_xer|out_data_buffer[14]~q ),
	.src_payload15(src_payload31),
	.out_data_buffer_15(\crosser_001|clock_xer|out_data_buffer[15]~q ),
	.src_payload16(src_payload32),
	.out_data_buffer_16(\crosser_001|clock_xer|out_data_buffer[16]~q ),
	.src_payload17(src_payload33),
	.out_data_buffer_17(\crosser_001|clock_xer|out_data_buffer[17]~q ),
	.src_payload18(src_payload34),
	.out_data_buffer_18(\crosser_001|clock_xer|out_data_buffer[18]~q ),
	.src_payload19(src_payload35),
	.out_data_buffer_19(\crosser_001|clock_xer|out_data_buffer[19]~q ),
	.src_payload20(src_payload36),
	.out_data_buffer_20(\crosser_001|clock_xer|out_data_buffer[20]~q ),
	.src_payload21(src_payload37),
	.out_data_buffer_21(\crosser_001|clock_xer|out_data_buffer[21]~q ),
	.src_payload22(src_payload38),
	.out_data_buffer_22(\crosser_001|clock_xer|out_data_buffer[22]~q ),
	.src_payload23(src_payload39),
	.out_data_buffer_23(\crosser_001|clock_xer|out_data_buffer[23]~q ),
	.src_payload24(src_payload40),
	.out_data_buffer_24(\crosser_001|clock_xer|out_data_buffer[24]~q ),
	.src_payload25(src_payload41),
	.out_data_buffer_25(\crosser_001|clock_xer|out_data_buffer[25]~q ),
	.src_payload26(src_payload42),
	.out_data_buffer_26(\crosser_001|clock_xer|out_data_buffer[26]~q ),
	.src_payload27(src_payload43),
	.out_data_buffer_27(\crosser_001|clock_xer|out_data_buffer[27]~q ),
	.src_payload28(src_payload44),
	.out_data_buffer_28(\crosser_001|clock_xer|out_data_buffer[28]~q ),
	.src_payload29(src_payload45),
	.out_data_buffer_29(\crosser_001|clock_xer|out_data_buffer[29]~q ),
	.src_payload30(src_payload46),
	.out_data_buffer_30(\crosser_001|clock_xer|out_data_buffer[30]~q ),
	.src_payload31(src_payload47),
	.out_data_buffer_31(\crosser_001|clock_xer|out_data_buffer[31]~q ),
	.src_payload32(src_payload48));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_4 cmd_mux_005(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.cp_valid(cp_valid),
	.F_pc_5(F_pc_5),
	.i_read(i_read),
	.read_accepted(\nios2_qsys_0_instruction_master_translator|read_accepted~q ),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.Equal0(Equal0),
	.rst1(rst1),
	.saved_grant_0(\cmd_mux_005|saved_grant[0]~q ),
	.mem_used_1(mem_used_15),
	.Equal1(\router_001|Equal1~1_combout ),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.WideOr11(WideOr13),
	.src_data_38(src_data_382),
	.src_data_39(src_data_392),
	.src4_valid(\cmd_demux_001|src4_valid~2_combout ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_3 cmd_mux_004(
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_31(d_writedata_31),
	.d_writedata_30(d_writedata_30),
	.d_writedata_29(d_writedata_29),
	.d_writedata_28(d_writedata_28),
	.d_writedata_27(d_writedata_27),
	.d_writedata_26(d_writedata_26),
	.d_writedata_25(d_writedata_25),
	.d_writedata_24(d_writedata_24),
	.cp_valid(cp_valid),
	.Equal8(\router|Equal8~4_combout ),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_3(F_pc_3),
	.F_pc_2(F_pc_2),
	.F_pc_4(F_pc_4),
	.d_writedata_0(d_writedata_0),
	.d_byteenable_0(d_byteenable_0),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.saved_grant_0(\cmd_mux_004|saved_grant[0]~q ),
	.waitrequest(waitrequest1),
	.mem_used_1(mem_used_14),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.src3_valid(\cmd_demux_001|src3_valid~0_combout ),
	.WideOr11(WideOr15),
	.hbreak_enabled(hbreak_enabled),
	.d_byteenable_2(d_byteenable_2),
	.src_data_46(src_data_461),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_21(d_writedata_21),
	.d_writedata_18(d_writedata_18),
	.d_writedata_23(d_writedata_23),
	.d_writedata_22(d_writedata_22),
	.d_writedata_20(d_writedata_20),
	.d_writedata_19(d_writedata_19),
	.src_payload(src_payload77),
	.src_payload1(src_payload78),
	.src_data_38(src_data_385),
	.src_data_39(src_data_395),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_32(src_data_322),
	.src_payload2(src_payload79),
	.src_payload3(src_payload80),
	.src_payload4(src_payload82),
	.src_payload5(src_payload83),
	.src_payload6(src_payload85),
	.src_data_33(src_data_331),
	.src_payload7(src_payload86),
	.src_payload8(src_payload87),
	.src_data_34(src_data_341),
	.src_payload9(src_payload88),
	.src_payload10(src_payload89),
	.src_payload11(src_payload90),
	.src_payload12(src_payload91),
	.src_payload13(src_payload92),
	.src_payload14(src_payload93),
	.src_payload15(src_payload94),
	.src_payload16(src_payload95),
	.src_data_35(src_data_351),
	.src_payload17(src_payload96),
	.src_payload18(src_payload97),
	.src_payload19(src_payload98),
	.src_payload20(src_payload99),
	.src_payload21(src_payload100),
	.src_payload22(src_payload101),
	.src_payload23(src_payload102),
	.src_payload24(src_payload103),
	.src_payload25(src_payload104),
	.src_payload26(src_payload105),
	.src_payload27(src_payload106),
	.src_payload28(src_payload107),
	.src_payload29(src_payload108),
	.src_payload30(src_payload109),
	.src_payload31(src_payload110),
	.src_payload32(src_payload111),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_2 cmd_mux_003(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_2(W_alu_result_2),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.F_pc_5(F_pc_5),
	.i_read(i_read),
	.read_accepted(\nios2_qsys_0_instruction_master_translator|read_accepted~q ),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.Equal0(Equal0),
	.uav_read1(uav_read),
	.rst1(rst1),
	.always1(\router|always1~0_combout ),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.Equal1(\router_001|Equal1~1_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.WideOr11(\cmd_mux_003|WideOr1~combout ),
	.wait_latency_counter_1(\sysid_qsys_0_control_slave_translator|wait_latency_counter[1]~0_combout ),
	.always11(\router_001|always1~1_combout ),
	.src_valid(\cmd_mux_003|src_valid~0_combout ),
	.src_data_68(\cmd_mux_003|src_data[68]~combout ),
	.always12(\router|always1~2_combout ),
	.src_payload(\cmd_mux_003|src_payload~0_combout ),
	.src_data_38(\cmd_mux_003|src_data[38]~combout ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_1 cmd_mux_001(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.saved_grant_1(saved_grant_1),
	.cp_valid(cp_valid),
	.Equal8(\router|Equal8~4_combout ),
	.Equal3(\router|Equal3~0_combout ),
	.Equal0(\router|Equal0~0_combout ),
	.src_valid(src_valid),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.src1_valid(src1_valid),
	.saved_grant_0(saved_grant_0),
	.mem_used_1(mem_used_1),
	.internal_reset(internal_reset),
	.d_byteenable_0(d_byteenable_0),
	.src_data_32(src_data_32),
	.F_pc_0(F_pc_0),
	.src_data_38(src_data_38),
	.F_pc_1(F_pc_1),
	.src_data_39(src_data_39),
	.r_sync_rst(r_sync_rst),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.WideOr11(WideOr1),
	.uav_read1(uav_read),
	.src_data_68(src_data_68),
	.waitrequest(waitrequest),
	.Equal2(Equal21),
	.s_serial_transferSTATE_1_PRE_WRITE(s_serial_transferSTATE_1_PRE_WRITE),
	.src_payload(src_payload6),
	.src_payload1(src_payload7),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux cmd_mux(
	.clk_0(clk_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.saved_grant_0(saved_grant_02),
	.out_data_buffer_3(out_data_buffer_3),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.out_data_buffer_38(\crosser_002|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_381(\crosser|clock_xer|out_data_buffer[38]~q ),
	.src_data_38(src_data_381),
	.out_data_buffer_39(\crosser_002|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_391(\crosser|clock_xer|out_data_buffer[39]~q ),
	.src_data_39(src_data_391),
	.out_valid(\crosser_002|clock_xer|out_valid~combout ),
	.out_data_toggle_flopped(\crosser|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid1(\crosser|clock_xer|out_valid~combout ),
	.WideOr11(WideOr12),
	.mem_used_1(mem_used_17),
	.last_cycle(last_cycle),
	.out_data_buffer_31(\crosser|clock_xer|out_data_buffer[31]~q ),
	.src_payload(src_payload5),
	.waitrequest_reset_override(\audio_avalon_audio_slave_translator|waitrequest_reset_override~q ),
	.out_data_buffer_107(\crosser_002|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_1071(\crosser|clock_xer|out_data_buffer[107]~q ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.out_data_buffer_68(\crosser_002|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_681(\crosser|clock_xer|out_data_buffer[68]~q ),
	.src_data_68(src_data_682),
	.out_data_buffer_30(\crosser|clock_xer|out_data_buffer[30]~q ),
	.src_payload1(src_payload16),
	.out_data_buffer_29(\crosser|clock_xer|out_data_buffer[29]~q ),
	.src_payload2(src_payload76),
	.out_data_buffer_28(\crosser|clock_xer|out_data_buffer[28]~q ),
	.src_payload3(src_payload81),
	.out_data_buffer_0(out_data_buffer_02),
	.out_data_buffer_1(out_data_buffer_110),
	.out_data_buffer_2(out_data_buffer_210),
	.out_data_buffer_27(\crosser|clock_xer|out_data_buffer[27]~q ),
	.src_payload4(src_payload84),
	.out_data_buffer_26(\crosser|clock_xer|out_data_buffer[26]~q ),
	.src_payload5(src_payload112),
	.out_data_buffer_25(\crosser|clock_xer|out_data_buffer[25]~q ),
	.src_payload6(src_payload113),
	.out_data_buffer_24(\crosser|clock_xer|out_data_buffer[24]~q ),
	.src_payload7(src_payload114),
	.out_data_buffer_23(\crosser|clock_xer|out_data_buffer[23]~q ),
	.src_payload8(src_payload115),
	.out_data_buffer_22(\crosser|clock_xer|out_data_buffer[22]~q ),
	.src_payload9(src_payload116),
	.out_data_buffer_21(\crosser|clock_xer|out_data_buffer[21]~q ),
	.src_payload10(src_payload117),
	.out_data_buffer_20(\crosser|clock_xer|out_data_buffer[20]~q ),
	.src_payload11(src_payload118),
	.out_data_buffer_19(\crosser|clock_xer|out_data_buffer[19]~q ),
	.src_payload12(src_payload119),
	.out_data_buffer_18(\crosser|clock_xer|out_data_buffer[18]~q ),
	.src_payload13(src_payload120),
	.out_data_buffer_17(\crosser|clock_xer|out_data_buffer[17]~q ),
	.src_payload14(src_payload121),
	.out_data_buffer_16(\crosser|clock_xer|out_data_buffer[16]~q ),
	.src_payload15(src_payload122),
	.out_data_buffer_15(\crosser|clock_xer|out_data_buffer[15]~q ),
	.src_payload16(src_payload123),
	.out_data_buffer_14(\crosser|clock_xer|out_data_buffer[14]~q ),
	.src_payload17(src_payload124),
	.out_data_buffer_13(\crosser|clock_xer|out_data_buffer[13]~q ),
	.src_payload18(src_payload125),
	.out_data_buffer_12(\crosser|clock_xer|out_data_buffer[12]~q ),
	.src_payload19(src_payload126),
	.out_data_buffer_11(\crosser|clock_xer|out_data_buffer[11]~q ),
	.src_payload20(src_payload127),
	.out_data_buffer_10(\crosser|clock_xer|out_data_buffer[10]~q ),
	.src_payload21(src_payload128),
	.out_data_buffer_9(\crosser|clock_xer|out_data_buffer[9]~q ),
	.src_payload22(src_payload129),
	.out_data_buffer_8(\crosser|clock_xer|out_data_buffer[8]~q ),
	.src_payload23(src_payload130),
	.out_data_buffer_7(\crosser|clock_xer|out_data_buffer[7]~q ),
	.src_payload24(src_payload131),
	.out_data_buffer_6(\crosser|clock_xer|out_data_buffer[6]~q ),
	.src_payload25(src_payload132),
	.out_data_buffer_5(\crosser|clock_xer|out_data_buffer[5]~q ),
	.src_payload26(src_payload133),
	.out_data_buffer_4(\crosser|clock_xer|out_data_buffer[4]~q ),
	.src_payload27(src_payload134),
	.src_payload28(src_payload135),
	.src_payload29(src_payload136),
	.src_payload30(src_payload137),
	.src_payload31(src_payload138));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.Equal5(\router_001|Equal5~4_combout ),
	.F_pc_10(F_pc_10),
	.Equal0(\router_001|Equal0~0_combout ),
	.F_pc_5(F_pc_5),
	.Equal01(\router_001|Equal0~1_combout ),
	.i_read(i_read),
	.read_accepted(\nios2_qsys_0_instruction_master_translator|read_accepted~q ),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.F_pc_2(F_pc_2),
	.F_pc_4(F_pc_4),
	.F_pc_9(F_pc_9),
	.src1_valid(src1_valid),
	.Equal1(\router_001|Equal1~1_combout ),
	.Equal02(\router_001|Equal0~3_combout ),
	.src_channel_6(\router_001|src_channel[6]~2_combout ),
	.Equal6(\router_001|Equal6~0_combout ),
	.src3_valid(\cmd_demux_001|src3_valid~0_combout ),
	.src6_valid(\cmd_demux_001|src6_valid~0_combout ),
	.src4_valid(\cmd_demux_001|src4_valid~2_combout ));

final_project_soc_final_project_soc_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.saved_grant_0(saved_grant_0),
	.uav_write(uav_write),
	.mem_used_1(mem_used_1),
	.Equal0(Equal0),
	.always0(always0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.always01(always01),
	.wait_latency_counter_11(wait_latency_counter_11),
	.wait_latency_counter_01(wait_latency_counter_01),
	.rst1(rst1),
	.always1(\router|always1~0_combout ),
	.Equal8(\router|Equal8~5_combout ),
	.src_channel_6(\router|src_channel[6]~7_combout ),
	.Equal01(\router|Equal0~3_combout ),
	.src_channel_9(\router|src_channel[9]~8_combout ),
	.in_ready(\crosser_001|clock_xer|in_ready~0_combout ),
	.WideOr0(\cmd_demux|WideOr0~2_combout ),
	.read_latency_shift_reg(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~2_combout ),
	.Equal3(\router|Equal3~1_combout ),
	.take_in_data(\crosser|clock_xer|take_in_data~0_combout ),
	.saved_grant_01(\cmd_mux_004|saved_grant[0]~q ),
	.waitrequest(waitrequest1),
	.mem_used_11(mem_used_14),
	.Equal1(\router|Equal1~0_combout ),
	.saved_grant_02(\cmd_mux_005|saved_grant[0]~q ),
	.mem_used_12(mem_used_15),
	.saved_grant_03(saved_grant_01),
	.mem_used_13(mem_used_16),
	.WideOr01(\cmd_demux|WideOr0~9_combout ),
	.saved_grant_04(\cmd_mux_003|saved_grant[0]~q ),
	.waitrequest1(waitrequest2),
	.cp_ready(\sysid_qsys_0_control_slave_agent|cp_ready~0_combout ),
	.WideOr02(\cmd_demux|WideOr0~10_combout ),
	.WideOr03(\cmd_demux|WideOr0~11_combout ));

final_project_soc_final_project_soc_mm_interconnect_0_router_002_5 router_008(
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.always0(\router_008|always0~0_combout ));

final_project_soc_final_project_soc_mm_interconnect_0_router_001 router_001(
	.F_pc_26(F_pc_26),
	.F_pc_25(F_pc_25),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.Equal5(\router_001|Equal5~4_combout ),
	.F_pc_10(F_pc_10),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.Equal0(\router_001|Equal0~0_combout ),
	.F_pc_5(F_pc_5),
	.F_pc_3(F_pc_3),
	.Equal01(\router_001|Equal0~1_combout ),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.F_pc_2(F_pc_2),
	.F_pc_4(F_pc_4),
	.F_pc_9(F_pc_9),
	.F_pc_1(F_pc_1),
	.Equal1(\router_001|Equal1~1_combout ),
	.always1(\router_001|always1~1_combout ),
	.Equal02(\router_001|Equal0~3_combout ),
	.src_channel_6(\router_001|src_channel[6]~2_combout ),
	.Equal6(\router_001|Equal6~0_combout ),
	.Equal2(\router_001|Equal2~1_combout ),
	.Equal51(\router_001|Equal5~5_combout ),
	.src_channel_5(\router_001|src_channel[5]~3_combout ));

final_project_soc_final_project_soc_mm_interconnect_0_router router(
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_3(W_alu_result_3),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.Equal8(\router|Equal8~4_combout ),
	.Equal3(\router|Equal3~0_combout ),
	.Equal0(\router|Equal0~0_combout ),
	.Equal01(Equal0),
	.Equal2(Equal2),
	.always1(\router|always1~0_combout ),
	.src_channel_6(\router|src_channel[6]~5_combout ),
	.src_channel_61(\router|src_channel[6]~6_combout ),
	.Equal81(\router|Equal8~5_combout ),
	.Equal21(\router|Equal2~3_combout ),
	.src_channel_62(\router|src_channel[6]~7_combout ),
	.Equal02(\router|Equal0~3_combout ),
	.src_channel_9(\router|src_channel[9]~8_combout ),
	.Equal22(Equal22),
	.Equal31(\router|Equal3~1_combout ),
	.Equal1(\router|Equal1~0_combout ),
	.always11(\router|always1~2_combout ));

final_project_soc_altera_avalon_sc_fifo_7 onchip_memory2_0_s1_agent_rsp_fifo(
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.uav_write(uav_write),
	.reset(r_sync_rst),
	.uav_read1(uav_read),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(mem_67_06),
	.rst1(rst1),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_16),
	.saved_grant_1(\cmd_mux_009|saved_grant[1]~q ),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ),
	.WideOr1(WideOr16),
	.mem1(\onchip_memory2_0_s1_agent_rsp_fifo|mem~1_combout ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_avalon_sc_fifo_4 ledg_s1_agent_rsp_fifo(
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.reset(r_sync_rst),
	.Equal0(Equal0),
	.mem_used_1(mem_used_11),
	.uav_read(uav_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.mem_67_0(mem_67_07),
	.rst1(rst1),
	.wait_latency_counter_0(\ledg_s1_translator|wait_latency_counter[0]~0_combout ),
	.read_latency_shift_reg(\ledg_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_avalon_sc_fifo_5 ledr_s1_agent_rsp_fifo(
	.W_alu_result_6(W_alu_result_6),
	.d_read(d_read),
	.d_write(d_write),
	.read_accepted(read_accepted),
	.write_accepted(write_accepted),
	.reset(r_sync_rst),
	.Equal2(Equal2),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.mem_67_0(mem_67_05),
	.rst1(rst1),
	.wait_latency_counter_0(\ledr_s1_translator|wait_latency_counter[0]~0_combout ),
	.read_latency_shift_reg(\ledr_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser_2 crosser_002(
	.clk_0(clk_0),
	.i_read(i_read),
	.read_accepted(\nios2_qsys_0_instruction_master_translator|read_accepted~q ),
	.F_pc_2(F_pc_2),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal2(\router_001|Equal2~1_combout ),
	.take_in_data(\crosser_002|clock_xer|take_in_data~2_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.out_data_buffer_38(\crosser_002|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser_002|clock_xer|out_data_buffer[39]~q ),
	.out_valid(\crosser_002|clock_xer|out_valid~combout ),
	.out_data_buffer_107(\crosser_002|clock_xer|out_data_buffer[107]~q ),
	.mem_used_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~0_combout ),
	.out_data_buffer_68(\crosser_002|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_86(\crosser_002|clock_xer|out_data_buffer[86]~q ),
	.clk_clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser_1 crosser_001(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.d_writedata_31(d_writedata_31),
	.d_writedata_30(d_writedata_30),
	.d_writedata_29(d_writedata_29),
	.d_writedata_28(d_writedata_28),
	.d_writedata_27(d_writedata_27),
	.d_writedata_26(d_writedata_26),
	.d_writedata_25(d_writedata_25),
	.d_writedata_24(d_writedata_24),
	.cp_valid(cp_valid),
	.uav_write(uav_write),
	.d_writedata_0(d_writedata_0),
	.d_byteenable_0(d_byteenable_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.uav_read(uav_read),
	.in_ready(\crosser_001|clock_xer|in_ready~0_combout ),
	.WideOr0(\cmd_demux|WideOr0~2_combout ),
	.last_cycle(last_cycle1),
	.saved_grant_0(\cmd_mux_006|saved_grant[0]~q ),
	.out_data_toggle_flopped(\crosser_001|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_001|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(\crosser_001|clock_xer|out_valid~combout ),
	.out_data_buffer_67(\crosser_001|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_68(\crosser_001|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_48(\crosser_001|clock_xer|out_data_buffer[48]~q ),
	.out_data_buffer_62(\crosser_001|clock_xer|out_data_buffer[62]~q ),
	.out_data_buffer_49(\crosser_001|clock_xer|out_data_buffer[49]~q ),
	.out_data_buffer_51(\crosser_001|clock_xer|out_data_buffer[51]~q ),
	.out_data_buffer_50(\crosser_001|clock_xer|out_data_buffer[50]~q ),
	.out_data_buffer_53(\crosser_001|clock_xer|out_data_buffer[53]~q ),
	.out_data_buffer_52(\crosser_001|clock_xer|out_data_buffer[52]~q ),
	.out_data_buffer_55(\crosser_001|clock_xer|out_data_buffer[55]~q ),
	.out_data_buffer_54(\crosser_001|clock_xer|out_data_buffer[54]~q ),
	.out_data_buffer_57(\crosser_001|clock_xer|out_data_buffer[57]~q ),
	.out_data_buffer_56(\crosser_001|clock_xer|out_data_buffer[56]~q ),
	.out_data_buffer_59(\crosser_001|clock_xer|out_data_buffer[59]~q ),
	.out_data_buffer_58(\crosser_001|clock_xer|out_data_buffer[58]~q ),
	.out_data_buffer_61(\crosser_001|clock_xer|out_data_buffer[61]~q ),
	.out_data_buffer_60(\crosser_001|clock_xer|out_data_buffer[60]~q ),
	.out_data_buffer_38(\crosser_001|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser_001|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_40(\crosser_001|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_41(\crosser_001|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_42(\crosser_001|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_43(\crosser_001|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_44(\crosser_001|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_45(\crosser_001|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_46(\crosser_001|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_47(\crosser_001|clock_xer|out_data_buffer[47]~q ),
	.out_data_buffer_32(out_data_buffer_32),
	.out_data_buffer_33(out_data_buffer_33),
	.out_data_buffer_34(out_data_buffer_34),
	.out_data_buffer_35(out_data_buffer_35),
	.out_data_buffer_107(\crosser_001|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_66(\crosser_001|clock_xer|out_data_buffer[66]~q ),
	.d_byteenable_2(d_byteenable_2),
	.WideOr01(\cmd_demux|WideOr0~11_combout ),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_3(d_byteenable_3),
	.out_data_buffer_0(\crosser_001|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser_001|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser_001|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser_001|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser_001|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser_001|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser_001|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser_001|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_8(\crosser_001|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_9(\crosser_001|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_10(\crosser_001|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_11(\crosser_001|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_12(\crosser_001|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_13(\crosser_001|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_14(\crosser_001|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_15(\crosser_001|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_16(\crosser_001|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_17(\crosser_001|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_18(\crosser_001|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_19(\crosser_001|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_20(\crosser_001|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_21(\crosser_001|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_22(\crosser_001|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_23(\crosser_001|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_24(\crosser_001|clock_xer|out_data_buffer[24]~q ),
	.out_data_buffer_25(\crosser_001|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_26(\crosser_001|clock_xer|out_data_buffer[26]~q ),
	.out_data_buffer_27(\crosser_001|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_28(\crosser_001|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_29(\crosser_001|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_30(\crosser_001|clock_xer|out_data_buffer[30]~q ),
	.out_data_buffer_31(\crosser_001|clock_xer|out_data_buffer[31]~q ),
	.d_writedata_21(d_writedata_21),
	.d_writedata_18(d_writedata_18),
	.d_writedata_23(d_writedata_23),
	.d_writedata_22(d_writedata_22),
	.d_writedata_20(d_writedata_20),
	.d_writedata_19(d_writedata_19),
	.clk_clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser crosser(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.clk_0(clk_0),
	.d_writedata_31(d_writedata_31),
	.d_writedata_30(d_writedata_30),
	.d_writedata_29(d_writedata_29),
	.d_writedata_28(d_writedata_28),
	.d_writedata_27(d_writedata_27),
	.d_writedata_26(d_writedata_26),
	.d_writedata_25(d_writedata_25),
	.d_writedata_24(d_writedata_24),
	.cp_valid(cp_valid),
	.uav_write(uav_write),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.uav_read(uav_read),
	.Equal3(\router|Equal3~1_combout ),
	.take_in_data(\crosser|clock_xer|take_in_data~0_combout ),
	.saved_grant_0(saved_grant_02),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_38(\crosser|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser|clock_xer|out_data_buffer[39]~q ),
	.out_data_toggle_flopped(\crosser|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(\crosser|clock_xer|out_valid~combout ),
	.out_data_buffer_67(\crosser|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_31(\crosser|clock_xer|out_data_buffer[31]~q ),
	.out_data_buffer_107(\crosser|clock_xer|out_data_buffer[107]~q ),
	.mem_used_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem_used[0]~0_combout ),
	.out_data_buffer_66(\crosser|clock_xer|out_data_buffer[66]~q ),
	.out_data_buffer_68(\crosser|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_30(\crosser|clock_xer|out_data_buffer[30]~q ),
	.d_writedata_21(d_writedata_21),
	.d_writedata_18(d_writedata_18),
	.d_writedata_23(d_writedata_23),
	.d_writedata_22(d_writedata_22),
	.d_writedata_20(d_writedata_20),
	.d_writedata_19(d_writedata_19),
	.out_data_buffer_29(\crosser|clock_xer|out_data_buffer[29]~q ),
	.out_data_buffer_28(\crosser|clock_xer|out_data_buffer[28]~q ),
	.out_data_buffer_0(out_data_buffer_02),
	.out_data_buffer_1(out_data_buffer_110),
	.out_data_buffer_2(out_data_buffer_210),
	.out_data_buffer_27(\crosser|clock_xer|out_data_buffer[27]~q ),
	.out_data_buffer_26(\crosser|clock_xer|out_data_buffer[26]~q ),
	.out_data_buffer_25(\crosser|clock_xer|out_data_buffer[25]~q ),
	.out_data_buffer_24(\crosser|clock_xer|out_data_buffer[24]~q ),
	.out_data_buffer_23(\crosser|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_22(\crosser|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_21(\crosser|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_20(\crosser|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_19(\crosser|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_18(\crosser|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_17(\crosser|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_16(\crosser|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_15(\crosser|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_14(\crosser|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_13(\crosser|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_12(\crosser|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_11(\crosser|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_10(\crosser|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_9(\crosser|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_8(\crosser|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_7(\crosser|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_6(\crosser|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_5(\crosser|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_4(\crosser|clock_xer|out_data_buffer[4]~q ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.readdata_16(readdata_16),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.read_latency_shift_reg_01(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_01(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_01(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.read_latency_shift_reg_02(read_latency_shift_reg_04),
	.mem_86_02(mem_86_01),
	.mem_68_02(mem_68_01),
	.src1_valid(src1_valid1),
	.src1_valid1(src1_valid2),
	.src1_valid2(src1_valid3),
	.src_payload(src_payload1),
	.src_payload1(src_payload2),
	.out_valid(out_valid2),
	.out_valid1(out_valid3),
	.WideOr11(\rsp_mux_001|WideOr1~combout ),
	.av_readdata_pre_30(av_readdata_pre_30),
	.src_payload2(src_payload4),
	.src_payload3(src_payload8),
	.readdata_5(readdata_51),
	.src_payload4(src_payload9));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_mux rsp_mux(
	.q_a_0(q_a_0),
	.readdata_0(readdata_0),
	.q_a_1(q_a_1),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.readdata_16(readdata_16),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.readdata_17(readdata_17),
	.q_a_17(q_a_17),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_23(q_a_23),
	.readdata_8(readdata_8),
	.q_a_8(q_a_8),
	.q_a_22(q_a_22),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.av_readdata_pre_16(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_22(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_20(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.src0_valid(src0_valid),
	.out_data_toggle_flopped(\crosser_004|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_004|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(out_valid),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_01(dreg_0),
	.out_valid1(out_valid1),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.read_latency_shift_reg_03(read_latency_shift_reg_03),
	.read_latency_shift_reg_04(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_01(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_01(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid1(src0_valid1),
	.src0_valid2(src0_valid2),
	.read_latency_shift_reg_05(read_latency_shift_reg_04),
	.mem_86_02(mem_86_01),
	.mem_68_02(mem_68_01),
	.src0_valid3(src0_valid3),
	.src0_valid4(src0_valid4),
	.WideOr11(WideOr11),
	.mem_67_0(mem_67_07),
	.src_payload(src_payload),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_01(av_readdata_pre_01),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.readdata_3(readdata_32),
	.av_readdata_pre_4(av_readdata_pre_4),
	.readdata_4(readdata_41),
	.av_readdata_pre_111(av_readdata_pre_111),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_161(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.readdata_5(readdata_51),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_211(av_readdata_pre_21),
	.av_readdata_pre_181(av_readdata_pre_18),
	.av_readdata_pre_171(av_readdata_pre_17),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_221(av_readdata_pre_22),
	.readdata_7(readdata_71),
	.av_readdata_pre_7(av_readdata_pre_7),
	.readdata_6(readdata_61),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_201(av_readdata_pre_20),
	.av_readdata_pre_191(av_readdata_pre_19),
	.src_payload1(src_payload10),
	.av_readdata_pre_02(\ledr_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.out_data_buffer_0(\crosser_006|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_01(\crosser_004|clock_xer|out_data_buffer[0]~q ),
	.av_readdata_pre_04(\ledg_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.src_data_1(src_data_1),
	.av_readdata_pre_110(\ledr_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_112(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_1(\crosser_006|clock_xer|out_data_buffer[1]~q ),
	.av_readdata_pre_113(\ledg_s1_translator|av_readdata_pre[1]~q ),
	.out_data_buffer_11(\crosser_004|clock_xer|out_data_buffer[1]~q ),
	.src_data_11(src_data_11),
	.src_data_2(src_data_2),
	.av_readdata_pre_24(\ledr_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_25(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_2(\crosser_006|clock_xer|out_data_buffer[2]~q ),
	.av_readdata_pre_26(\ledg_s1_translator|av_readdata_pre[2]~q ),
	.out_data_buffer_21(\crosser_004|clock_xer|out_data_buffer[2]~q ),
	.src_data_21(src_data_21),
	.src_data_3(src_data_3),
	.av_readdata_pre_31(\ledr_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_3(\crosser_006|clock_xer|out_data_buffer[3]~q ),
	.av_readdata_pre_33(\ledg_s1_translator|av_readdata_pre[3]~q ),
	.out_data_buffer_31(\crosser_004|clock_xer|out_data_buffer[3]~q ),
	.src_data_31(src_data_31),
	.src_data_4(src_data_4),
	.av_readdata_pre_41(\ledr_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_42(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.out_data_buffer_4(\crosser_006|clock_xer|out_data_buffer[4]~q ),
	.av_readdata_pre_43(\ledg_s1_translator|av_readdata_pre[4]~q ),
	.out_data_buffer_41(\crosser_004|clock_xer|out_data_buffer[4]~q ),
	.src_data_41(src_data_410),
	.av_readdata_pre_51(\ledr_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.out_data_buffer_5(\crosser_006|clock_xer|out_data_buffer[5]~q ),
	.av_readdata_pre_53(\ledg_s1_translator|av_readdata_pre[5]~q ),
	.out_data_buffer_51(\crosser_004|clock_xer|out_data_buffer[5]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_61(\ledr_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_6(\crosser_006|clock_xer|out_data_buffer[6]~q ),
	.av_readdata_pre_63(\ledg_s1_translator|av_readdata_pre[6]~q ),
	.out_data_buffer_61(\crosser_004|clock_xer|out_data_buffer[6]~q ),
	.src_data_61(src_data_63),
	.av_readdata_pre_71(\ledr_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_72(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.out_data_buffer_7(\crosser_006|clock_xer|out_data_buffer[7]~q ),
	.av_readdata_pre_73(\ledg_s1_translator|av_readdata_pre[7]~q ),
	.out_data_buffer_71(\crosser_004|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_8(\crosser_004|clock_xer|out_data_buffer[8]~q ),
	.av_readdata_pre_81(\ledr_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.out_data_buffer_81(\crosser_006|clock_xer|out_data_buffer[8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_91(\ledr_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.out_data_buffer_9(\crosser_006|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_91(\crosser_004|clock_xer|out_data_buffer[9]~q ),
	.src_data_9(src_data_9),
	.out_data_buffer_10(\crosser_004|clock_xer|out_data_buffer[10]~q ),
	.av_readdata_pre_101(\ledr_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_102(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.out_data_buffer_101(\crosser_006|clock_xer|out_data_buffer[10]~q ),
	.src_data_10(src_data_10),
	.out_data_buffer_111(\crosser_006|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_112(\crosser_004|clock_xer|out_data_buffer[11]~q ),
	.av_readdata_pre_114(\ledr_s1_translator|av_readdata_pre[11]~q ),
	.src_data_111(src_data_111),
	.av_readdata_pre_121(\ledr_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_122(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.out_data_buffer_12(\crosser_006|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_121(\crosser_004|clock_xer|out_data_buffer[12]~q ),
	.src_data_12(src_data_12),
	.av_readdata_pre_131(\ledr_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_132(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.out_data_buffer_13(\crosser_006|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_131(\crosser_004|clock_xer|out_data_buffer[13]~q ),
	.src_data_13(src_data_13),
	.out_data_buffer_14(\crosser_004|clock_xer|out_data_buffer[14]~q ),
	.av_readdata_pre_141(\ledr_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_142(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.out_data_buffer_141(\crosser_006|clock_xer|out_data_buffer[14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_151(\ledr_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_152(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.out_data_buffer_15(\crosser_006|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_151(\crosser_004|clock_xer|out_data_buffer[15]~q ),
	.src_data_15(src_data_15),
	.out_data_buffer_16(\crosser_004|clock_xer|out_data_buffer[16]~q ),
	.av_readdata_pre_162(\ledr_s1_translator|av_readdata_pre[16]~q ),
	.out_data_buffer_161(\crosser_006|clock_xer|out_data_buffer[16]~q ),
	.src_data_16(src_data_16),
	.out_data_buffer_17(\crosser_004|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_171(\crosser_006|clock_xer|out_data_buffer[17]~q ),
	.av_readdata_pre_172(\ledr_s1_translator|av_readdata_pre[17]~q ),
	.src_data_17(src_data_17),
	.out_data_buffer_23(\crosser_004|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_231(\crosser_006|clock_xer|out_data_buffer[23]~q ),
	.src_data_23(src_data_23),
	.out_data_buffer_22(\crosser_004|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_221(\crosser_006|clock_xer|out_data_buffer[22]~q ),
	.src_data_22(src_data_22),
	.out_data_buffer_211(\crosser_006|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_212(\crosser_004|clock_xer|out_data_buffer[21]~q ),
	.src_data_211(src_data_211),
	.out_data_buffer_20(\crosser_006|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_201(\crosser_004|clock_xer|out_data_buffer[20]~q ),
	.src_data_20(src_data_20),
	.out_data_buffer_19(\crosser_006|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_191(\crosser_004|clock_xer|out_data_buffer[19]~q ),
	.src_data_19(src_data_19),
	.out_data_buffer_18(\crosser_004|clock_xer|out_data_buffer[18]~q ),
	.out_data_buffer_181(\crosser_006|clock_xer|out_data_buffer[18]~q ),
	.src_data_18(src_data_18),
	.src_data_51(src_data_510),
	.src_data_71(src_data_71));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_5 rsp_demux_009(
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid4),
	.src1_valid(src1_valid3));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_4 rsp_demux_006(
	.mem_86_0(\sdram_s1_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sdram_s1_agent_rsp_fifo|mem[0][68]~q ),
	.in_data_toggle(\crosser_007|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_007|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.in_data_toggle1(\crosser_006|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_006|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.always0(\router_008|always0~0_combout ),
	.WideOr0(\rsp_demux_006|WideOr0~1_combout ));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_3 rsp_demux_005(
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.mem_86_0(mem_86_01),
	.mem_68_0(mem_68_01),
	.src0_valid(src0_valid3));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_2 rsp_demux_004(
	.read_latency_shift_reg_0(\nios2_qsys_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\nios2_qsys_0_debug_mem_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid2),
	.src1_valid(src1_valid2));

final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_1 rsp_demux_003(
	.read_latency_shift_reg_0(\sysid_qsys_0_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_86_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\sysid_qsys_0_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(src0_valid1));

final_project_soc_altera_avalon_st_handshake_clock_crosser_7 crosser_007(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.out_valid(out_valid3),
	.out_data_buffer_67(\crosser_007|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_11),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_36),
	.out_data_buffer_4(out_data_buffer_41),
	.in_data_toggle(\crosser_007|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_007|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.always0(\router_008|always0~0_combout ),
	.mem_67_0(\sdram_s1_agent_rsp_fifo|mem[0][67]~q ),
	.take_in_data(\crosser_006|clock_xer|take_in_data~0_combout ),
	.out_data_buffer_11(out_data_buffer_111),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_141),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_21(out_data_buffer_211),
	.out_data_buffer_18(out_data_buffer_181),
	.out_data_buffer_17(out_data_buffer_171),
	.out_data_buffer_31(out_data_buffer_311),
	.out_data_buffer_30(out_data_buffer_301),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_28(out_data_buffer_281),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_261),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_10(out_data_buffer_101),
	.out_data_buffer_24(out_data_buffer_241),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_8(out_data_buffer_81),
	.out_data_buffer_22(out_data_buffer_221),
	.out_data_buffer_7(out_data_buffer_71),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_payload_0(\sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.out_payload_1(\sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.out_payload_2(\sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.out_payload_3(\sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.out_payload_4(\sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.out_payload_11(\sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.out_payload_13(\sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.out_payload_16(\sdram_s1_agent_rdata_fifo|out_payload[16]~q ),
	.out_payload_12(\sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.out_payload_5(\sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.out_payload_14(\sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.out_payload_15(\sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.out_payload_21(\sdram_s1_agent_rdata_fifo|out_payload[21]~q ),
	.out_payload_18(\sdram_s1_agent_rdata_fifo|out_payload[18]~q ),
	.out_payload_17(\sdram_s1_agent_rdata_fifo|out_payload[17]~q ),
	.out_payload_31(\sdram_s1_agent_rdata_fifo|out_payload[31]~q ),
	.out_payload_30(\sdram_s1_agent_rdata_fifo|out_payload[30]~q ),
	.out_payload_29(\sdram_s1_agent_rdata_fifo|out_payload[29]~q ),
	.out_payload_28(\sdram_s1_agent_rdata_fifo|out_payload[28]~q ),
	.out_payload_27(\sdram_s1_agent_rdata_fifo|out_payload[27]~q ),
	.out_payload_26(\sdram_s1_agent_rdata_fifo|out_payload[26]~q ),
	.out_payload_25(\sdram_s1_agent_rdata_fifo|out_payload[25]~q ),
	.out_payload_10(\sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.out_payload_24(\sdram_s1_agent_rdata_fifo|out_payload[24]~q ),
	.out_payload_9(\sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.out_payload_23(\sdram_s1_agent_rdata_fifo|out_payload[23]~q ),
	.out_payload_8(\sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.out_payload_22(\sdram_s1_agent_rdata_fifo|out_payload[22]~q ),
	.out_payload_7(\sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.out_payload_6(\sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.out_payload_20(\sdram_s1_agent_rdata_fifo|out_payload[20]~q ),
	.out_payload_19(\sdram_s1_agent_rdata_fifo|out_payload[19]~q ),
	.clk_clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser_6 crosser_006(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid(out_valid1),
	.out_data_buffer_67(out_data_buffer_671),
	.mem_used_0(\sdram_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_107_0(\sdram_s1_agent_rsp_fifo|mem[0][107]~q ),
	.out_valid1(\sdram_s1_agent_rdata_fifo|out_valid~q ),
	.in_data_toggle(\crosser_006|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_006|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.always0(\router_008|always0~0_combout ),
	.mem_67_0(\sdram_s1_agent_rsp_fifo|mem[0][67]~q ),
	.take_in_data(\crosser_006|clock_xer|take_in_data~0_combout ),
	.out_data_buffer_0(\crosser_006|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser_006|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser_006|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser_006|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser_006|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser_006|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser_006|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser_006|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_8(\crosser_006|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_9(\crosser_006|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_10(\crosser_006|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_11(\crosser_006|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_12(\crosser_006|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_13(\crosser_006|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_14(\crosser_006|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_15(\crosser_006|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_16(\crosser_006|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_17(\crosser_006|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_28(out_data_buffer_282),
	.out_data_buffer_27(out_data_buffer_272),
	.out_data_buffer_26(out_data_buffer_262),
	.out_data_buffer_25(out_data_buffer_252),
	.out_data_buffer_24(out_data_buffer_242),
	.out_data_buffer_23(\crosser_006|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_22(\crosser_006|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_21(\crosser_006|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_20(\crosser_006|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_19(\crosser_006|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_18(\crosser_006|clock_xer|out_data_buffer[18]~q ),
	.out_payload_0(\sdram_s1_agent_rdata_fifo|out_payload[0]~q ),
	.out_payload_1(\sdram_s1_agent_rdata_fifo|out_payload[1]~q ),
	.out_payload_2(\sdram_s1_agent_rdata_fifo|out_payload[2]~q ),
	.out_payload_3(\sdram_s1_agent_rdata_fifo|out_payload[3]~q ),
	.out_payload_4(\sdram_s1_agent_rdata_fifo|out_payload[4]~q ),
	.out_payload_11(\sdram_s1_agent_rdata_fifo|out_payload[11]~q ),
	.out_payload_13(\sdram_s1_agent_rdata_fifo|out_payload[13]~q ),
	.out_payload_16(\sdram_s1_agent_rdata_fifo|out_payload[16]~q ),
	.out_payload_12(\sdram_s1_agent_rdata_fifo|out_payload[12]~q ),
	.out_payload_5(\sdram_s1_agent_rdata_fifo|out_payload[5]~q ),
	.out_payload_14(\sdram_s1_agent_rdata_fifo|out_payload[14]~q ),
	.out_payload_15(\sdram_s1_agent_rdata_fifo|out_payload[15]~q ),
	.out_payload_21(\sdram_s1_agent_rdata_fifo|out_payload[21]~q ),
	.out_payload_18(\sdram_s1_agent_rdata_fifo|out_payload[18]~q ),
	.out_payload_17(\sdram_s1_agent_rdata_fifo|out_payload[17]~q ),
	.out_payload_31(\sdram_s1_agent_rdata_fifo|out_payload[31]~q ),
	.out_payload_30(\sdram_s1_agent_rdata_fifo|out_payload[30]~q ),
	.out_payload_29(\sdram_s1_agent_rdata_fifo|out_payload[29]~q ),
	.out_payload_28(\sdram_s1_agent_rdata_fifo|out_payload[28]~q ),
	.out_data_buffer_31(out_data_buffer_313),
	.out_payload_27(\sdram_s1_agent_rdata_fifo|out_payload[27]~q ),
	.out_data_buffer_30(out_data_buffer_302),
	.out_payload_26(\sdram_s1_agent_rdata_fifo|out_payload[26]~q ),
	.out_data_buffer_29(out_data_buffer_292),
	.out_payload_25(\sdram_s1_agent_rdata_fifo|out_payload[25]~q ),
	.out_payload_10(\sdram_s1_agent_rdata_fifo|out_payload[10]~q ),
	.out_payload_24(\sdram_s1_agent_rdata_fifo|out_payload[24]~q ),
	.out_payload_9(\sdram_s1_agent_rdata_fifo|out_payload[9]~q ),
	.out_payload_23(\sdram_s1_agent_rdata_fifo|out_payload[23]~q ),
	.out_payload_8(\sdram_s1_agent_rdata_fifo|out_payload[8]~q ),
	.out_payload_22(\sdram_s1_agent_rdata_fifo|out_payload[22]~q ),
	.out_payload_7(\sdram_s1_agent_rdata_fifo|out_payload[7]~q ),
	.out_payload_6(\sdram_s1_agent_rdata_fifo|out_payload[6]~q ),
	.out_payload_20(\sdram_s1_agent_rdata_fifo|out_payload[20]~q ),
	.out_payload_19(\sdram_s1_agent_rdata_fifo|out_payload[19]~q ),
	.clk_clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser_5 crosser_005(
	.clk_0(clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid2),
	.out_data_buffer_67(\crosser_005|clock_xer|out_data_buffer[67]~q ),
	.out_data_buffer_0(out_data_buffer_01),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_21),
	.out_data_buffer_3(out_data_buffer_31),
	.out_data_buffer_4(out_data_buffer_4),
	.mem_86_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][86]~q ),
	.mem_68_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][68]~q ),
	.in_data_toggle(\crosser_005|clock_xer|in_data_toggle~q ),
	.dreg_0(\crosser_005|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.take_in_data(\crosser_005|clock_xer|take_in_data~0_combout ),
	.mem_67_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][67]~q ),
	.rp_valid(\audio_avalon_audio_slave_agent|rp_valid~combout ),
	.out_data_buffer_11(out_data_buffer_112),
	.out_data_buffer_13(out_data_buffer_131),
	.out_data_buffer_16(out_data_buffer_161),
	.out_data_buffer_12(out_data_buffer_121),
	.out_data_buffer_5(out_data_buffer_51),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_151),
	.out_data_buffer_21(out_data_buffer_212),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_31(out_data_buffer_312),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_291),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_271),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_251),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_9(out_data_buffer_91),
	.out_data_buffer_23(out_data_buffer_231),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_61),
	.out_data_buffer_20(out_data_buffer_201),
	.out_data_buffer_19(out_data_buffer_191),
	.out_data_0(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_11(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[11]~5_combout ),
	.out_data_13(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[13]~6_combout ),
	.out_data_16(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[16]~7_combout ),
	.out_data_12(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[12]~8_combout ),
	.out_data_5(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[5]~9_combout ),
	.out_data_14(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[14]~10_combout ),
	.out_data_15(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[15]~11_combout ),
	.out_data_21(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[21]~12_combout ),
	.out_data_18(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[18]~13_combout ),
	.out_data_17(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[17]~14_combout ),
	.out_data_31(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[31]~15_combout ),
	.out_data_30(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[30]~16_combout ),
	.out_data_29(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[29]~17_combout ),
	.out_data_28(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[28]~18_combout ),
	.out_data_27(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[27]~19_combout ),
	.out_data_26(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[26]~20_combout ),
	.out_data_25(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[25]~21_combout ),
	.out_data_10(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[10]~22_combout ),
	.out_data_24(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[24]~23_combout ),
	.out_data_9(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[9]~24_combout ),
	.out_data_23(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[23]~25_combout ),
	.out_data_8(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[8]~26_combout ),
	.out_data_22(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[22]~27_combout ),
	.out_data_7(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[7]~28_combout ),
	.out_data_6(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[6]~29_combout ),
	.out_data_20(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[20]~30_combout ),
	.out_data_19(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[19]~31_combout ),
	.clk_clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser_4 crosser_004(
	.clk_0(clk_0),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped(\crosser_004|clock_xer|out_data_toggle_flopped~q ),
	.dreg_0(\crosser_004|clock_xer|in_to_out_synchronizer|dreg[0]~q ),
	.out_valid(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.in_data_toggle(\crosser_004|clock_xer|in_data_toggle~q ),
	.dreg_01(\crosser_004|clock_xer|out_to_in_synchronizer|dreg[0]~q ),
	.take_in_data(\crosser_005|clock_xer|take_in_data~0_combout ),
	.mem_67_0(\audio_avalon_audio_slave_agent_rsp_fifo|mem[0][67]~q ),
	.rp_valid(\audio_avalon_audio_slave_agent|rp_valid~combout ),
	.out_data_buffer_0(\crosser_004|clock_xer|out_data_buffer[0]~q ),
	.out_data_buffer_1(\crosser_004|clock_xer|out_data_buffer[1]~q ),
	.out_data_buffer_2(\crosser_004|clock_xer|out_data_buffer[2]~q ),
	.out_data_buffer_3(\crosser_004|clock_xer|out_data_buffer[3]~q ),
	.out_data_buffer_4(\crosser_004|clock_xer|out_data_buffer[4]~q ),
	.out_data_buffer_5(\crosser_004|clock_xer|out_data_buffer[5]~q ),
	.out_data_buffer_6(\crosser_004|clock_xer|out_data_buffer[6]~q ),
	.out_data_buffer_7(\crosser_004|clock_xer|out_data_buffer[7]~q ),
	.out_data_buffer_8(\crosser_004|clock_xer|out_data_buffer[8]~q ),
	.out_data_buffer_9(\crosser_004|clock_xer|out_data_buffer[9]~q ),
	.out_data_buffer_10(\crosser_004|clock_xer|out_data_buffer[10]~q ),
	.out_data_buffer_11(\crosser_004|clock_xer|out_data_buffer[11]~q ),
	.out_data_buffer_12(\crosser_004|clock_xer|out_data_buffer[12]~q ),
	.out_data_buffer_13(\crosser_004|clock_xer|out_data_buffer[13]~q ),
	.out_data_buffer_14(\crosser_004|clock_xer|out_data_buffer[14]~q ),
	.out_data_buffer_15(\crosser_004|clock_xer|out_data_buffer[15]~q ),
	.out_data_buffer_16(\crosser_004|clock_xer|out_data_buffer[16]~q ),
	.out_data_buffer_17(\crosser_004|clock_xer|out_data_buffer[17]~q ),
	.out_data_buffer_28(out_data_buffer_283),
	.out_data_buffer_27(out_data_buffer_273),
	.out_data_buffer_26(out_data_buffer_263),
	.out_data_buffer_25(out_data_buffer_253),
	.out_data_buffer_24(out_data_buffer_243),
	.out_data_buffer_23(\crosser_004|clock_xer|out_data_buffer[23]~q ),
	.out_data_buffer_22(\crosser_004|clock_xer|out_data_buffer[22]~q ),
	.out_data_buffer_21(\crosser_004|clock_xer|out_data_buffer[21]~q ),
	.out_data_buffer_20(\crosser_004|clock_xer|out_data_buffer[20]~q ),
	.out_data_buffer_19(\crosser_004|clock_xer|out_data_buffer[19]~q ),
	.out_data_buffer_18(\crosser_004|clock_xer|out_data_buffer[18]~q ),
	.out_data_0(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_11(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[11]~5_combout ),
	.out_data_13(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[13]~6_combout ),
	.out_data_16(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[16]~7_combout ),
	.out_data_12(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[12]~8_combout ),
	.out_data_5(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[5]~9_combout ),
	.out_data_14(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[14]~10_combout ),
	.out_data_15(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[15]~11_combout ),
	.out_data_21(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[21]~12_combout ),
	.out_data_18(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[18]~13_combout ),
	.out_data_17(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[17]~14_combout ),
	.out_data_31(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[31]~15_combout ),
	.out_data_30(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[30]~16_combout ),
	.out_data_29(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[29]~17_combout ),
	.out_data_28(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[28]~18_combout ),
	.out_data_buffer_31(out_data_buffer_314),
	.out_data_27(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[27]~19_combout ),
	.out_data_buffer_30(out_data_buffer_303),
	.out_data_26(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[26]~20_combout ),
	.out_data_buffer_29(out_data_buffer_293),
	.out_data_25(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[25]~21_combout ),
	.out_data_10(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[10]~22_combout ),
	.out_data_24(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[24]~23_combout ),
	.out_data_9(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[9]~24_combout ),
	.out_data_23(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[23]~25_combout ),
	.out_data_8(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[8]~26_combout ),
	.out_data_22(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[22]~27_combout ),
	.out_data_7(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[7]~28_combout ),
	.out_data_6(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[6]~29_combout ),
	.out_data_20(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[20]~30_combout ),
	.out_data_19(\audio_avalon_audio_slave_agent_rdata_fifo|out_data[19]~31_combout ),
	.clk_clk(clk_clk));

final_project_soc_altera_avalon_st_handshake_clock_crosser_3 crosser_003(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_3(F_pc_3),
	.uav_read(\nios2_qsys_0_instruction_master_translator|uav_read~combout ),
	.F_pc_2(F_pc_2),
	.F_pc_4(F_pc_4),
	.F_pc_9(F_pc_9),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.src_channel_5(\router_001|src_channel[5]~3_combout ),
	.in_ready(\crosser_003|clock_xer|in_ready~0_combout ),
	.last_cycle(last_cycle1),
	.saved_grant_1(saved_grant_11),
	.out_valid(\crosser_003|clock_xer|out_valid~combout ),
	.out_data_buffer_68(\crosser_003|clock_xer|out_data_buffer[68]~q ),
	.out_data_buffer_48(\crosser_003|clock_xer|out_data_buffer[48]~q ),
	.out_data_buffer_62(\crosser_003|clock_xer|out_data_buffer[62]~q ),
	.out_data_buffer_49(\crosser_003|clock_xer|out_data_buffer[49]~q ),
	.out_data_buffer_51(\crosser_003|clock_xer|out_data_buffer[51]~q ),
	.out_data_buffer_50(\crosser_003|clock_xer|out_data_buffer[50]~q ),
	.out_data_buffer_53(\crosser_003|clock_xer|out_data_buffer[53]~q ),
	.out_data_buffer_52(\crosser_003|clock_xer|out_data_buffer[52]~q ),
	.out_data_buffer_55(\crosser_003|clock_xer|out_data_buffer[55]~q ),
	.out_data_buffer_54(\crosser_003|clock_xer|out_data_buffer[54]~q ),
	.out_data_buffer_57(\crosser_003|clock_xer|out_data_buffer[57]~q ),
	.out_data_buffer_56(\crosser_003|clock_xer|out_data_buffer[56]~q ),
	.out_data_buffer_59(\crosser_003|clock_xer|out_data_buffer[59]~q ),
	.out_data_buffer_58(\crosser_003|clock_xer|out_data_buffer[58]~q ),
	.out_data_buffer_61(\crosser_003|clock_xer|out_data_buffer[61]~q ),
	.out_data_buffer_60(\crosser_003|clock_xer|out_data_buffer[60]~q ),
	.out_data_buffer_38(\crosser_003|clock_xer|out_data_buffer[38]~q ),
	.out_data_buffer_39(\crosser_003|clock_xer|out_data_buffer[39]~q ),
	.out_data_buffer_40(\crosser_003|clock_xer|out_data_buffer[40]~q ),
	.out_data_buffer_41(\crosser_003|clock_xer|out_data_buffer[41]~q ),
	.out_data_buffer_42(\crosser_003|clock_xer|out_data_buffer[42]~q ),
	.out_data_buffer_43(\crosser_003|clock_xer|out_data_buffer[43]~q ),
	.out_data_buffer_44(\crosser_003|clock_xer|out_data_buffer[44]~q ),
	.out_data_buffer_45(\crosser_003|clock_xer|out_data_buffer[45]~q ),
	.out_data_buffer_46(\crosser_003|clock_xer|out_data_buffer[46]~q ),
	.out_data_buffer_47(\crosser_003|clock_xer|out_data_buffer[47]~q ),
	.out_data_buffer_32(out_data_buffer_321),
	.out_data_buffer_33(out_data_buffer_331),
	.out_data_buffer_34(out_data_buffer_341),
	.out_data_buffer_35(out_data_buffer_351),
	.out_data_buffer_107(\crosser_003|clock_xer|out_data_buffer[107]~q ),
	.out_data_buffer_86(\crosser_003|clock_xer|out_data_buffer[86]~q ),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_sc_fifo (
	clk,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_21,
	readdata_18,
	readdata_17,
	readdata_31,
	readdata_30,
	readdata_29,
	readdata_28,
	readdata_27,
	readdata_26,
	readdata_25,
	readdata_10,
	readdata_24,
	readdata_9,
	readdata_23,
	readdata_8,
	readdata_22,
	readdata_7,
	readdata_6,
	readdata_20,
	readdata_19,
	reset,
	mem_used_0,
	mem_107_0,
	read_latency_shift_reg_0,
	mem_used_01,
	rp_valid,
	WideOr0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_11,
	out_data_13,
	out_data_16,
	out_data_12,
	out_data_5,
	out_data_14,
	out_data_15,
	out_data_21,
	out_data_18,
	out_data_17,
	out_data_31,
	out_data_30,
	out_data_29,
	out_data_28,
	out_data_27,
	out_data_26,
	out_data_25,
	out_data_10,
	out_data_24,
	out_data_9,
	out_data_23,
	out_data_8,
	out_data_22,
	out_data_7,
	out_data_6,
	out_data_20,
	out_data_19)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	readdata_0;
input 	readdata_1;
input 	readdata_2;
input 	readdata_3;
input 	readdata_4;
input 	readdata_11;
input 	readdata_13;
input 	readdata_16;
input 	readdata_12;
input 	readdata_5;
input 	readdata_14;
input 	readdata_15;
input 	readdata_21;
input 	readdata_18;
input 	readdata_17;
input 	readdata_31;
input 	readdata_30;
input 	readdata_29;
input 	readdata_28;
input 	readdata_27;
input 	readdata_26;
input 	readdata_25;
input 	readdata_10;
input 	readdata_24;
input 	readdata_9;
input 	readdata_23;
input 	readdata_8;
input 	readdata_22;
input 	readdata_7;
input 	readdata_6;
input 	readdata_20;
input 	readdata_19;
input 	reset;
input 	mem_used_0;
input 	mem_107_0;
input 	read_latency_shift_reg_0;
output 	mem_used_01;
input 	rp_valid;
input 	WideOr0;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_11;
output 	out_data_13;
output 	out_data_16;
output 	out_data_12;
output 	out_data_5;
output 	out_data_14;
output 	out_data_15;
output 	out_data_21;
output 	out_data_18;
output 	out_data_17;
output 	out_data_31;
output 	out_data_30;
output 	out_data_29;
output 	out_data_28;
output 	out_data_27;
output 	out_data_26;
output 	out_data_25;
output 	out_data_10;
output 	out_data_24;
output 	out_data_9;
output 	out_data_23;
output 	out_data_8;
output 	out_data_22;
output 	out_data_7;
output 	out_data_6;
output 	out_data_20;
output 	out_data_19;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[0][0]~q ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[0][1]~q ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[0][2]~q ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[0][3]~q ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[0][4]~q ;
wire \mem[1][11]~q ;
wire \mem~5_combout ;
wire \mem[0][11]~q ;
wire \mem[1][13]~q ;
wire \mem~6_combout ;
wire \mem[0][13]~q ;
wire \mem[1][16]~q ;
wire \mem~7_combout ;
wire \mem[0][16]~q ;
wire \mem[1][12]~q ;
wire \mem~8_combout ;
wire \mem[0][12]~q ;
wire \mem[1][5]~q ;
wire \mem~9_combout ;
wire \mem[0][5]~q ;
wire \mem[1][14]~q ;
wire \mem~10_combout ;
wire \mem[0][14]~q ;
wire \mem[1][15]~q ;
wire \mem~11_combout ;
wire \mem[0][15]~q ;
wire \mem[1][21]~q ;
wire \mem~12_combout ;
wire \mem[0][21]~q ;
wire \mem[1][18]~q ;
wire \mem~13_combout ;
wire \mem[0][18]~q ;
wire \mem[1][17]~q ;
wire \mem~14_combout ;
wire \mem[0][17]~q ;
wire \mem[1][31]~q ;
wire \mem~15_combout ;
wire \mem[0][31]~q ;
wire \mem[1][30]~q ;
wire \mem~16_combout ;
wire \mem[0][30]~q ;
wire \mem[1][29]~q ;
wire \mem~17_combout ;
wire \mem[0][29]~q ;
wire \mem[1][28]~q ;
wire \mem~18_combout ;
wire \mem[0][28]~q ;
wire \mem[1][27]~q ;
wire \mem~19_combout ;
wire \mem[0][27]~q ;
wire \mem[1][26]~q ;
wire \mem~20_combout ;
wire \mem[0][26]~q ;
wire \mem[1][25]~q ;
wire \mem~21_combout ;
wire \mem[0][25]~q ;
wire \mem[1][10]~q ;
wire \mem~22_combout ;
wire \mem[0][10]~q ;
wire \mem[1][24]~q ;
wire \mem~23_combout ;
wire \mem[0][24]~q ;
wire \mem[1][9]~q ;
wire \mem~24_combout ;
wire \mem[0][9]~q ;
wire \mem[1][23]~q ;
wire \mem~25_combout ;
wire \mem[0][23]~q ;
wire \mem[1][8]~q ;
wire \mem~26_combout ;
wire \mem[0][8]~q ;
wire \mem[1][22]~q ;
wire \mem~27_combout ;
wire \mem[0][22]~q ;
wire \mem[1][7]~q ;
wire \mem~28_combout ;
wire \mem[0][7]~q ;
wire \mem[1][6]~q ;
wire \mem~29_combout ;
wire \mem[0][6]~q ;
wire \mem[1][20]~q ;
wire \mem~30_combout ;
wire \mem[0][20]~q ;
wire \mem[1][19]~q ;
wire \mem~31_combout ;
wire \mem[0][19]~q ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_01),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \out_data[0]~0 (
	.dataa(\mem[0][0]~q ),
	.datab(readdata_0),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0]~0 .lut_mask = 16'hEFFE;
defparam \out_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[1]~1 (
	.dataa(\mem[0][1]~q ),
	.datab(readdata_1),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1]~1 .lut_mask = 16'hEFFE;
defparam \out_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[2]~2 (
	.dataa(\mem[0][2]~q ),
	.datab(readdata_2),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_2),
	.cout());
defparam \out_data[2]~2 .lut_mask = 16'hEFFE;
defparam \out_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[3]~3 (
	.dataa(\mem[0][3]~q ),
	.datab(readdata_3),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_3),
	.cout());
defparam \out_data[3]~3 .lut_mask = 16'hEFFE;
defparam \out_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[4]~4 (
	.dataa(\mem[0][4]~q ),
	.datab(readdata_4),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_4),
	.cout());
defparam \out_data[4]~4 .lut_mask = 16'hEFFE;
defparam \out_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[11]~5 (
	.dataa(\mem[0][11]~q ),
	.datab(readdata_11),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_11),
	.cout());
defparam \out_data[11]~5 .lut_mask = 16'hEFFE;
defparam \out_data[11]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[13]~6 (
	.dataa(\mem[0][13]~q ),
	.datab(readdata_13),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_13),
	.cout());
defparam \out_data[13]~6 .lut_mask = 16'hEFFE;
defparam \out_data[13]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[16]~7 (
	.dataa(\mem[0][16]~q ),
	.datab(readdata_16),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_16),
	.cout());
defparam \out_data[16]~7 .lut_mask = 16'hEFFE;
defparam \out_data[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[12]~8 (
	.dataa(\mem[0][12]~q ),
	.datab(readdata_12),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_12),
	.cout());
defparam \out_data[12]~8 .lut_mask = 16'hEFFE;
defparam \out_data[12]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[5]~9 (
	.dataa(\mem[0][5]~q ),
	.datab(readdata_5),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5]~9 .lut_mask = 16'hEFFE;
defparam \out_data[5]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[14]~10 (
	.dataa(\mem[0][14]~q ),
	.datab(readdata_14),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_14),
	.cout());
defparam \out_data[14]~10 .lut_mask = 16'hEFFE;
defparam \out_data[14]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[15]~11 (
	.dataa(\mem[0][15]~q ),
	.datab(readdata_15),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_15),
	.cout());
defparam \out_data[15]~11 .lut_mask = 16'hEFFE;
defparam \out_data[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[21]~12 (
	.dataa(\mem[0][21]~q ),
	.datab(readdata_21),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_21),
	.cout());
defparam \out_data[21]~12 .lut_mask = 16'hEFFE;
defparam \out_data[21]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[18]~13 (
	.dataa(\mem[0][18]~q ),
	.datab(readdata_18),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_18),
	.cout());
defparam \out_data[18]~13 .lut_mask = 16'hEFFE;
defparam \out_data[18]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[17]~14 (
	.dataa(\mem[0][17]~q ),
	.datab(readdata_17),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_17),
	.cout());
defparam \out_data[17]~14 .lut_mask = 16'hEFFE;
defparam \out_data[17]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[31]~15 (
	.dataa(\mem[0][31]~q ),
	.datab(readdata_31),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_31),
	.cout());
defparam \out_data[31]~15 .lut_mask = 16'hEFFE;
defparam \out_data[31]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[30]~16 (
	.dataa(\mem[0][30]~q ),
	.datab(readdata_30),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_30),
	.cout());
defparam \out_data[30]~16 .lut_mask = 16'hEFFE;
defparam \out_data[30]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[29]~17 (
	.dataa(\mem[0][29]~q ),
	.datab(readdata_29),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_29),
	.cout());
defparam \out_data[29]~17 .lut_mask = 16'hEFFE;
defparam \out_data[29]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[28]~18 (
	.dataa(\mem[0][28]~q ),
	.datab(readdata_28),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_28),
	.cout());
defparam \out_data[28]~18 .lut_mask = 16'hEFFE;
defparam \out_data[28]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[27]~19 (
	.dataa(\mem[0][27]~q ),
	.datab(readdata_27),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_27),
	.cout());
defparam \out_data[27]~19 .lut_mask = 16'hEFFE;
defparam \out_data[27]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[26]~20 (
	.dataa(\mem[0][26]~q ),
	.datab(readdata_26),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_26),
	.cout());
defparam \out_data[26]~20 .lut_mask = 16'hEFFE;
defparam \out_data[26]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[25]~21 (
	.dataa(\mem[0][25]~q ),
	.datab(readdata_25),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_25),
	.cout());
defparam \out_data[25]~21 .lut_mask = 16'hEFFE;
defparam \out_data[25]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[10]~22 (
	.dataa(\mem[0][10]~q ),
	.datab(readdata_10),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_10),
	.cout());
defparam \out_data[10]~22 .lut_mask = 16'hEFFE;
defparam \out_data[10]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[24]~23 (
	.dataa(\mem[0][24]~q ),
	.datab(readdata_24),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_24),
	.cout());
defparam \out_data[24]~23 .lut_mask = 16'hEFFE;
defparam \out_data[24]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[9]~24 (
	.dataa(\mem[0][9]~q ),
	.datab(readdata_9),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_9),
	.cout());
defparam \out_data[9]~24 .lut_mask = 16'hEFFE;
defparam \out_data[9]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[23]~25 (
	.dataa(\mem[0][23]~q ),
	.datab(readdata_23),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_23),
	.cout());
defparam \out_data[23]~25 .lut_mask = 16'hEFFE;
defparam \out_data[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[8]~26 (
	.dataa(\mem[0][8]~q ),
	.datab(readdata_8),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_8),
	.cout());
defparam \out_data[8]~26 .lut_mask = 16'hEFFE;
defparam \out_data[8]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[22]~27 (
	.dataa(\mem[0][22]~q ),
	.datab(readdata_22),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_22),
	.cout());
defparam \out_data[22]~27 .lut_mask = 16'hEFFE;
defparam \out_data[22]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[7]~28 (
	.dataa(\mem[0][7]~q ),
	.datab(readdata_7),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_7),
	.cout());
defparam \out_data[7]~28 .lut_mask = 16'hEFFE;
defparam \out_data[7]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[6]~29 (
	.dataa(\mem[0][6]~q ),
	.datab(readdata_6),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_6),
	.cout());
defparam \out_data[6]~29 .lut_mask = 16'hEFFE;
defparam \out_data[6]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[20]~30 (
	.dataa(\mem[0][20]~q ),
	.datab(readdata_20),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_20),
	.cout());
defparam \out_data[20]~30 .lut_mask = 16'hEFFE;
defparam \out_data[20]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[19]~31 (
	.dataa(\mem[0][19]~q ),
	.datab(readdata_19),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(out_data_19),
	.cout());
defparam \out_data[19]~31 .lut_mask = 16'hEFFE;
defparam \out_data[19]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(mem_used_0),
	.datab(mem_107_0),
	.datac(WideOr0),
	.datad(rp_valid),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h7FFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~q ),
	.datab(read_latency_shift_reg_0),
	.datac(mem_used_01),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~0 (
	.dataa(\mem_used[1]~q ),
	.datab(mem_used_01),
	.datac(read_latency_shift_reg_0),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~0_combout ),
	.cout());
defparam \mem_used[0]~0 .lut_mask = 16'hFDFE;
defparam \mem_used[0]~0 .sum_lutc_input = "datac";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][0]~q ),
	.datab(readdata_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][1]~q ),
	.datab(readdata_1),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][2]~q ),
	.datab(readdata_2),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][2]~q ),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][3]~q ),
	.datab(readdata_3),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][3]~q ),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][4]~q ),
	.datab(readdata_4),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][4]~q ),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[1][11]~q ),
	.datab(readdata_11),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hAACC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][11]~q ),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[1][13]~q ),
	.datab(readdata_13),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][13]~q ),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[1][16]~q ),
	.datab(readdata_16),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hAACC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][16]~q ),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[1][12]~q ),
	.datab(readdata_12),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hAACC;
defparam \mem~8 .sum_lutc_input = "datac";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][12]~q ),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[1][5]~q ),
	.datab(readdata_5),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hAACC;
defparam \mem~9 .sum_lutc_input = "datac";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][5]~q ),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[1][14]~q ),
	.datab(readdata_14),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hAACC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][14]~q ),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[1][15]~q ),
	.datab(readdata_15),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hAACC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][15]~q ),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[1][21]~q ),
	.datab(readdata_21),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][21]~q ),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[1][18]~q ),
	.datab(readdata_18),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hAACC;
defparam \mem~13 .sum_lutc_input = "datac";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][18]~q ),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[1][17]~q ),
	.datab(readdata_17),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][17]~q ),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[1][31]~q ),
	.datab(readdata_31),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hAACC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][31]~q ),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[1][30]~q ),
	.datab(readdata_30),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAACC;
defparam \mem~16 .sum_lutc_input = "datac";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][30]~q ),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[1][29]~q ),
	.datab(readdata_29),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hAACC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][29]~q ),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[1][28]~q ),
	.datab(readdata_28),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][28]~q ),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[1][27]~q ),
	.datab(readdata_27),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hAACC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][27]~q ),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[1][26]~q ),
	.datab(readdata_26),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][26]~q ),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[1][25]~q ),
	.datab(readdata_25),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hAACC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][25]~q ),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cycloneive_lcell_comb \mem~22 (
	.dataa(\mem[1][10]~q ),
	.datab(readdata_10),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~22_combout ),
	.cout());
defparam \mem~22 .lut_mask = 16'hAACC;
defparam \mem~22 .sum_lutc_input = "datac";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][10]~q ),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cycloneive_lcell_comb \mem~23 (
	.dataa(\mem[1][24]~q ),
	.datab(readdata_24),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~23_combout ),
	.cout());
defparam \mem~23 .lut_mask = 16'hAACC;
defparam \mem~23 .sum_lutc_input = "datac";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][24]~q ),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cycloneive_lcell_comb \mem~24 (
	.dataa(\mem[1][9]~q ),
	.datab(readdata_9),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~24_combout ),
	.cout());
defparam \mem~24 .lut_mask = 16'hAACC;
defparam \mem~24 .sum_lutc_input = "datac";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][9]~q ),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cycloneive_lcell_comb \mem~25 (
	.dataa(\mem[1][23]~q ),
	.datab(readdata_23),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~25_combout ),
	.cout());
defparam \mem~25 .lut_mask = 16'hAACC;
defparam \mem~25 .sum_lutc_input = "datac";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][23]~q ),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cycloneive_lcell_comb \mem~26 (
	.dataa(\mem[1][8]~q ),
	.datab(readdata_8),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~26_combout ),
	.cout());
defparam \mem~26 .lut_mask = 16'hAACC;
defparam \mem~26 .sum_lutc_input = "datac";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][8]~q ),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cycloneive_lcell_comb \mem~27 (
	.dataa(\mem[1][22]~q ),
	.datab(readdata_22),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~27_combout ),
	.cout());
defparam \mem~27 .lut_mask = 16'hAACC;
defparam \mem~27 .sum_lutc_input = "datac";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][22]~q ),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cycloneive_lcell_comb \mem~28 (
	.dataa(\mem[1][7]~q ),
	.datab(readdata_7),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~28_combout ),
	.cout());
defparam \mem~28 .lut_mask = 16'hAACC;
defparam \mem~28 .sum_lutc_input = "datac";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][7]~q ),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cycloneive_lcell_comb \mem~29 (
	.dataa(\mem[1][6]~q ),
	.datab(readdata_6),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~29_combout ),
	.cout());
defparam \mem~29 .lut_mask = 16'hAACC;
defparam \mem~29 .sum_lutc_input = "datac";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][6]~q ),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cycloneive_lcell_comb \mem~30 (
	.dataa(\mem[1][20]~q ),
	.datab(readdata_20),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~30_combout ),
	.cout());
defparam \mem~30 .lut_mask = 16'hAACC;
defparam \mem~30 .sum_lutc_input = "datac";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][20]~q ),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cycloneive_lcell_comb \mem~31 (
	.dataa(\mem[1][19]~q ),
	.datab(readdata_19),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~31_combout ),
	.cout());
defparam \mem~31 .lut_mask = 16'hAACC;
defparam \mem~31 .sum_lutc_input = "datac";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][19]~q ),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

endmodule

module final_project_soc_altera_avalon_sc_fifo_1 (
	clk,
	reset,
	saved_grant_0,
	saved_grant_1,
	WideOr1,
	mem_used_1,
	out_data_buffer_67,
	waitrequest_reset_override,
	mem_used_0,
	mem_used_01,
	mem_107_0,
	rp_valid,
	mem_86_0,
	mem_68_0,
	WideOr0,
	sink_ready,
	nonposted_write_endofpacket,
	src_data_68,
	mem_67_0,
	out_data_buffer_86)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	saved_grant_0;
input 	saved_grant_1;
input 	WideOr1;
output 	mem_used_1;
input 	out_data_buffer_67;
input 	waitrequest_reset_override;
output 	mem_used_0;
output 	mem_used_01;
output 	mem_107_0;
input 	rp_valid;
output 	mem_86_0;
output 	mem_68_0;
input 	WideOr0;
input 	sink_ready;
input 	nonposted_write_endofpacket;
input 	src_data_68;
output 	mem_67_0;
input 	out_data_buffer_86;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[1]~3_combout ;
wire \mem_used[1]~4_combout ;
wire \mem_used[0]~5_combout ;
wire \mem_used[0]~6_combout ;
wire \mem[1][107]~q ;
wire \mem~0_combout ;
wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;
wire \mem[1][67]~q ;
wire \mem~3_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~0 (
	.dataa(waitrequest_reset_override),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(mem_used_0),
	.cout());
defparam \mem_used[0]~0 .lut_mask = 16'hAAFF;
defparam \mem_used[0]~0 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_01),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~3_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~3_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~3_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~3_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(mem_used_01),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(nonposted_write_endofpacket),
	.datab(WideOr1),
	.datac(src_data_68),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFE;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~3 (
	.dataa(mem_used_01),
	.datab(WideOr0),
	.datac(rp_valid),
	.datad(mem_107_0),
	.cin(gnd),
	.combout(\mem_used[1]~3_combout ),
	.cout());
defparam \mem_used[1]~3 .lut_mask = 16'hFF7F;
defparam \mem_used[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~4 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(waitrequest_reset_override),
	.datac(\mem_used[0]~2_combout ),
	.datad(\mem_used[1]~3_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~4_combout ),
	.cout());
defparam \mem_used[1]~4 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~5 (
	.dataa(mem_used_0),
	.datab(nonposted_write_endofpacket),
	.datac(WideOr1),
	.datad(src_data_68),
	.cin(gnd),
	.combout(\mem_used[0]~5_combout ),
	.cout());
defparam \mem_used[0]~5 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~6 (
	.dataa(\mem_used[0]~5_combout ),
	.datab(mem_used_01),
	.datac(mem_used_1),
	.datad(sink_ready),
	.cin(gnd),
	.combout(\mem_used[0]~6_combout ),
	.cout());
defparam \mem_used[0]~6 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~6 .sum_lutc_input = "datac";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hFAFC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFAFC;
defparam \mem~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_2 (
	saved_grant_1,
	saved_grant_0,
	uav_write,
	mem_used_1,
	reset,
	WideOr1,
	src_data_68,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	waitrequest,
	clk)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_1;
input 	saved_grant_0;
input 	uav_write;
output 	mem_used_1;
input 	reset;
input 	WideOr1;
input 	src_data_68;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	waitrequest;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][86]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~2_combout ;
wire \mem[1][68]~q ;
wire \mem~1_combout ;
wire \mem[1][67]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~2_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~2_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~2_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(WideOr1),
	.datab(src_data_68),
	.datac(waitrequest),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEFEF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~3_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hBF8F;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(src_data_68),
	.datab(WideOr1),
	.datac(waitrequest),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hEFEF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hFF55;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][67]~q ),
	.datab(saved_grant_0),
	.datac(uav_write),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hFAFC;
defparam \mem~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_3 (
	d_read,
	d_write,
	read_accepted,
	write_accepted,
	reset,
	uav_read,
	read_latency_shift_reg_0,
	mem_67_0,
	Equal2,
	av_waitrequest,
	mem_used_1,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	d_write;
input 	read_accepted;
input 	write_accepted;
input 	reset;
input 	uav_read;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	Equal2;
input 	av_waitrequest;
output 	mem_used_1;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem[1][67]~q ;
wire \mem~2_combout ;
wire \mem[0][67]~3_combout ;
wire \mem_used[1]~4_combout ;
wire \mem_used[1]~5_combout ;


dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(d_read),
	.datab(read_accepted),
	.datac(\mem_used[0]~2_combout ),
	.datad(read_latency_shift_reg),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFFFB;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hB8FF;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(read_latency_shift_reg_0),
	.datac(mem_67_0),
	.datad(\mem~2_combout ),
	.cin(gnd),
	.combout(\mem[0][67]~3_combout ),
	.cout());
defparam \mem[0][67]~3 .lut_mask = 16'hFFF6;
defparam \mem[0][67]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~4 (
	.dataa(\mem_used[0]~q ),
	.datab(av_waitrequest),
	.datac(Equal2),
	.datad(uav_read),
	.cin(gnd),
	.combout(\mem_used[1]~4_combout ),
	.cout());
defparam \mem_used[1]~4 .lut_mask = 16'hFFFD;
defparam \mem_used[1]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~5 (
	.dataa(\mem_used[0]~q ),
	.datab(\mem_used[1]~4_combout ),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[1]~5_combout ),
	.cout());
defparam \mem_used[1]~5 .lut_mask = 16'hDF8F;
defparam \mem_used[1]~5 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_4 (
	W_alu_result_7,
	W_alu_result_5,
	d_write,
	write_accepted,
	reset,
	Equal0,
	mem_used_1,
	uav_read,
	read_latency_shift_reg_0,
	mem_67_0,
	rst1,
	wait_latency_counter_0,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	d_write;
input 	write_accepted;
input 	reset;
input 	Equal0;
output 	mem_used_1;
input 	uav_read;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	rst1;
input 	wait_latency_counter_0;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem[1][67]~q ;
wire \mem~0_combout ;
wire \mem[0][67]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(W_alu_result_7),
	.datab(W_alu_result_5),
	.datac(rst1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFBFB;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(Equal0),
	.datab(uav_read),
	.datac(wait_latency_counter_0),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFFFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~1_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hB8FF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_5 (
	W_alu_result_6,
	d_read,
	d_write,
	read_accepted,
	write_accepted,
	reset,
	Equal2,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_67_0,
	rst1,
	wait_latency_counter_0,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_6;
input 	d_read;
input 	d_write;
input 	read_accepted;
input 	write_accepted;
input 	reset;
input 	Equal2;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_67_0;
input 	rst1;
input 	wait_latency_counter_0;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~5_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~3_combout ;
wire \mem[1][67]~q ;
wire \mem~0_combout ;
wire \mem[0][67]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem[0][67]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~5 (
	.dataa(d_read),
	.datab(read_accepted),
	.datac(W_alu_result_6),
	.datad(rst1),
	.cin(gnd),
	.combout(\mem_used[1]~5_combout ),
	.cout());
defparam \mem_used[1]~5 .lut_mask = 16'hFFFB;
defparam \mem_used[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(Equal2),
	.datab(wait_latency_counter_0),
	.datac(\mem_used[1]~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hFEFE;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~3 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~2_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~3_combout ),
	.cout());
defparam \mem_used[1]~3 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~3 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][67]~q ),
	.datab(mem_used_1),
	.datac(d_write),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hB8FF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem[0][67]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_67_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][67]~1_combout ),
	.cout());
defparam \mem[0][67]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][67]~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_6 (
	d_write,
	write_accepted,
	uav_read,
	uav_write,
	reset,
	uav_read1,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_1,
	mem,
	local_read,
	mem1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	uav_read;
input 	uav_write;
input 	reset;
input 	uav_read1;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
input 	saved_grant_1;
output 	mem;
input 	local_read;
output 	mem1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;
wire \mem[1][67]~q ;
wire \mem~3_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hFFFE;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~4 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(write_accepted),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(mem1),
	.cout());
defparam \mem~4 .lut_mask = 16'hEFFF;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(local_read),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hEFFF;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][68]~q ),
	.datab(mem),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFAFC;
defparam \mem~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(local_read),
	.datac(\mem_used[1]~0_combout ),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_7 (
	uav_read,
	uav_write,
	reset,
	uav_read1,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	rst1,
	saved_grant_0,
	mem_used_1,
	saved_grant_1,
	mem,
	WideOr1,
	mem1,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	uav_read;
input 	uav_write;
input 	reset;
input 	uav_read1;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	rst1;
input 	saved_grant_0;
output 	mem_used_1;
input 	saved_grant_1;
output 	mem;
input 	WideOr1;
output 	mem1;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~3_combout ;
wire \mem[1][67]~q ;
wire \mem~4_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(saved_grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hAAFF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~1 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(mem1),
	.cout());
defparam \mem~1 .lut_mask = 16'hFFFE;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][68]~q ),
	.datab(mem1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hFAFC;
defparam \mem~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(mem1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~1_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_8 (
	d_write,
	write_accepted,
	uav_read,
	uav_write,
	reset,
	uav_read1,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	rst1,
	saved_grant_0,
	mem_used_1,
	saved_grant_1,
	WideOr1,
	mem,
	mem1,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	uav_read;
input 	uav_write;
input 	reset;
input 	uav_read1;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	rst1;
input 	saved_grant_0;
output 	mem_used_1;
input 	saved_grant_1;
input 	WideOr1;
output 	mem;
output 	mem1;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~3_combout ;
wire \mem[1][67]~q ;
wire \mem~4_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(write_accepted),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~0 .lut_mask = 16'hEFFF;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~1 (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(mem1),
	.cout());
defparam \mem~1 .lut_mask = 16'hFFFE;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][68]~q ),
	.datab(mem1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hFAFC;
defparam \mem~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(mem1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hFEFE;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~1_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_9 (
	clk,
	reset,
	mem_used_0,
	mem_107_0,
	out_valid1,
	WideOr0,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_11,
	out_payload_13,
	out_payload_16,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_21,
	out_payload_18,
	out_payload_17,
	out_payload_31,
	out_payload_30,
	out_payload_29,
	out_payload_28,
	out_payload_27,
	out_payload_26,
	out_payload_25,
	out_payload_10,
	out_payload_24,
	out_payload_9,
	out_payload_23,
	out_payload_8,
	out_payload_22,
	out_payload_7,
	out_payload_6,
	out_payload_20,
	out_payload_19,
	za_valid,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_11,
	za_data_13,
	za_data_16,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_21,
	za_data_18,
	za_data_17,
	za_data_31,
	za_data_30,
	za_data_29,
	za_data_28,
	za_data_27,
	za_data_26,
	za_data_25,
	za_data_10,
	za_data_24,
	za_data_9,
	za_data_23,
	za_data_8,
	za_data_22,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_19)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	mem_used_0;
input 	mem_107_0;
output 	out_valid1;
input 	WideOr0;
output 	out_payload_0;
output 	out_payload_1;
output 	out_payload_2;
output 	out_payload_3;
output 	out_payload_4;
output 	out_payload_11;
output 	out_payload_13;
output 	out_payload_16;
output 	out_payload_12;
output 	out_payload_5;
output 	out_payload_14;
output 	out_payload_15;
output 	out_payload_21;
output 	out_payload_18;
output 	out_payload_17;
output 	out_payload_31;
output 	out_payload_30;
output 	out_payload_29;
output 	out_payload_28;
output 	out_payload_27;
output 	out_payload_26;
output 	out_payload_25;
output 	out_payload_10;
output 	out_payload_24;
output 	out_payload_9;
output 	out_payload_23;
output 	out_payload_8;
output 	out_payload_22;
output 	out_payload_7;
output 	out_payload_6;
output 	out_payload_20;
output 	out_payload_19;
input 	za_valid;
input 	za_data_0;
input 	za_data_1;
input 	za_data_2;
input 	za_data_3;
input 	za_data_4;
input 	za_data_11;
input 	za_data_13;
input 	za_data_16;
input 	za_data_12;
input 	za_data_5;
input 	za_data_14;
input 	za_data_15;
input 	za_data_21;
input 	za_data_18;
input 	za_data_17;
input 	za_data_31;
input 	za_data_30;
input 	za_data_29;
input 	za_data_28;
input 	za_data_27;
input 	za_data_26;
input 	za_data_25;
input 	za_data_10;
input 	za_data_24;
input 	za_data_9;
input 	za_data_23;
input 	za_data_8;
input 	za_data_22;
input 	za_data_7;
input 	za_data_6;
input 	za_data_20;
input 	za_data_19;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \internal_out_ready~0_combout ;
wire \mem_rd_ptr[0]~1_combout ;
wire \rd_ptr[0]~q ;
wire \mem_rd_ptr[1]~0_combout ;
wire \rd_ptr[1]~q ;
wire \wr_ptr[0]~0_combout ;
wire \next_full~0_combout ;
wire \read~0_combout ;
wire \mem_rd_ptr[2]~2_combout ;
wire \rd_ptr[2]~q ;
wire \wr_ptr[2]~q ;
wire \Add0~1_combout ;
wire \next_full~1_combout ;
wire \next_full~2_combout ;
wire \full~q ;
wire \write~combout ;
wire \wr_ptr[0]~q ;
wire \Add0~0_combout ;
wire \wr_ptr[1]~q ;
wire \internal_out_valid~0_combout ;
wire \Equal0~0_combout ;
wire \internal_out_valid~1_combout ;
wire \next_empty~0_combout ;
wire \empty~q ;
wire \internal_out_valid~2_combout ;
wire \internal_out_valid~q ;
wire \mem~416_combout ;
wire \mem~160_q ;
wire \mem~417_combout ;
wire \mem~192_q ;
wire \mem~418_combout ;
wire \mem~128_q ;
wire \mem~256_combout ;
wire \mem~419_combout ;
wire \mem~224_q ;
wire \mem~257_combout ;
wire \mem~420_combout ;
wire \mem~64_q ;
wire \mem~421_combout ;
wire \mem~32_q ;
wire \mem~422_combout ;
wire \mem~0_q ;
wire \mem~258_combout ;
wire \mem~423_combout ;
wire \mem~96_q ;
wire \mem~259_combout ;
wire \mem~260_combout ;
wire \internal_out_payload[0]~q ;
wire \mem~161_q ;
wire \mem~193_q ;
wire \mem~129_q ;
wire \mem~261_combout ;
wire \mem~225_q ;
wire \mem~262_combout ;
wire \mem~65_q ;
wire \mem~33_q ;
wire \mem~1_q ;
wire \mem~263_combout ;
wire \mem~97_q ;
wire \mem~264_combout ;
wire \mem~265_combout ;
wire \internal_out_payload[1]~q ;
wire \mem~162_q ;
wire \mem~194_q ;
wire \mem~130_q ;
wire \mem~266_combout ;
wire \mem~226_q ;
wire \mem~267_combout ;
wire \mem~66_q ;
wire \mem~34_q ;
wire \mem~2_q ;
wire \mem~268_combout ;
wire \mem~98_q ;
wire \mem~269_combout ;
wire \mem~270_combout ;
wire \internal_out_payload[2]~q ;
wire \mem~163_q ;
wire \mem~195_q ;
wire \mem~131_q ;
wire \mem~271_combout ;
wire \mem~227_q ;
wire \mem~272_combout ;
wire \mem~67_q ;
wire \mem~35_q ;
wire \mem~3_q ;
wire \mem~273_combout ;
wire \mem~99_q ;
wire \mem~274_combout ;
wire \mem~275_combout ;
wire \internal_out_payload[3]~q ;
wire \mem~164_q ;
wire \mem~196_q ;
wire \mem~132_q ;
wire \mem~276_combout ;
wire \mem~228_q ;
wire \mem~277_combout ;
wire \mem~68_q ;
wire \mem~36_q ;
wire \mem~4_q ;
wire \mem~278_combout ;
wire \mem~100_q ;
wire \mem~279_combout ;
wire \mem~280_combout ;
wire \internal_out_payload[4]~q ;
wire \mem~171_q ;
wire \mem~203_q ;
wire \mem~139_q ;
wire \mem~281_combout ;
wire \mem~235_q ;
wire \mem~282_combout ;
wire \mem~75_q ;
wire \mem~43_q ;
wire \mem~11_q ;
wire \mem~283_combout ;
wire \mem~107_q ;
wire \mem~284_combout ;
wire \mem~285_combout ;
wire \internal_out_payload[11]~q ;
wire \mem~173_q ;
wire \mem~205_q ;
wire \mem~141_q ;
wire \mem~286_combout ;
wire \mem~237_q ;
wire \mem~287_combout ;
wire \mem~77_q ;
wire \mem~45_q ;
wire \mem~13_q ;
wire \mem~288_combout ;
wire \mem~109_q ;
wire \mem~289_combout ;
wire \mem~290_combout ;
wire \internal_out_payload[13]~q ;
wire \mem~176_q ;
wire \mem~208_q ;
wire \mem~144_q ;
wire \mem~291_combout ;
wire \mem~240_q ;
wire \mem~292_combout ;
wire \mem~80_q ;
wire \mem~48_q ;
wire \mem~16_q ;
wire \mem~293_combout ;
wire \mem~112_q ;
wire \mem~294_combout ;
wire \mem~295_combout ;
wire \internal_out_payload[16]~q ;
wire \mem~172_q ;
wire \mem~204_q ;
wire \mem~140_q ;
wire \mem~296_combout ;
wire \mem~236_q ;
wire \mem~297_combout ;
wire \mem~76_q ;
wire \mem~44_q ;
wire \mem~12_q ;
wire \mem~298_combout ;
wire \mem~108_q ;
wire \mem~299_combout ;
wire \mem~300_combout ;
wire \internal_out_payload[12]~q ;
wire \mem~165_q ;
wire \mem~197_q ;
wire \mem~133_q ;
wire \mem~301_combout ;
wire \mem~229_q ;
wire \mem~302_combout ;
wire \mem~69_q ;
wire \mem~37_q ;
wire \mem~5_q ;
wire \mem~303_combout ;
wire \mem~101_q ;
wire \mem~304_combout ;
wire \mem~305_combout ;
wire \internal_out_payload[5]~q ;
wire \mem~174_q ;
wire \mem~206_q ;
wire \mem~142_q ;
wire \mem~306_combout ;
wire \mem~238_q ;
wire \mem~307_combout ;
wire \mem~78_q ;
wire \mem~46_q ;
wire \mem~14_q ;
wire \mem~308_combout ;
wire \mem~110_q ;
wire \mem~309_combout ;
wire \mem~310_combout ;
wire \internal_out_payload[14]~q ;
wire \mem~175_q ;
wire \mem~207_q ;
wire \mem~143_q ;
wire \mem~311_combout ;
wire \mem~239_q ;
wire \mem~312_combout ;
wire \mem~79_q ;
wire \mem~47_q ;
wire \mem~15_q ;
wire \mem~313_combout ;
wire \mem~111_q ;
wire \mem~314_combout ;
wire \mem~315_combout ;
wire \internal_out_payload[15]~q ;
wire \mem~181_q ;
wire \mem~213_q ;
wire \mem~149_q ;
wire \mem~316_combout ;
wire \mem~245_q ;
wire \mem~317_combout ;
wire \mem~85_q ;
wire \mem~53_q ;
wire \mem~21_q ;
wire \mem~318_combout ;
wire \mem~117_q ;
wire \mem~319_combout ;
wire \mem~320_combout ;
wire \internal_out_payload[21]~q ;
wire \mem~178_q ;
wire \mem~210_q ;
wire \mem~146_q ;
wire \mem~321_combout ;
wire \mem~242_q ;
wire \mem~322_combout ;
wire \mem~82_q ;
wire \mem~50_q ;
wire \mem~18_q ;
wire \mem~323_combout ;
wire \mem~114_q ;
wire \mem~324_combout ;
wire \mem~325_combout ;
wire \internal_out_payload[18]~q ;
wire \mem~177_q ;
wire \mem~209_q ;
wire \mem~145_q ;
wire \mem~326_combout ;
wire \mem~241_q ;
wire \mem~327_combout ;
wire \mem~81_q ;
wire \mem~49_q ;
wire \mem~17_q ;
wire \mem~328_combout ;
wire \mem~113_q ;
wire \mem~329_combout ;
wire \mem~330_combout ;
wire \internal_out_payload[17]~q ;
wire \mem~191_q ;
wire \mem~223_q ;
wire \mem~159_q ;
wire \mem~331_combout ;
wire \mem~255_q ;
wire \mem~332_combout ;
wire \mem~95_q ;
wire \mem~63_q ;
wire \mem~31_q ;
wire \mem~333_combout ;
wire \mem~127_q ;
wire \mem~334_combout ;
wire \mem~335_combout ;
wire \internal_out_payload[31]~q ;
wire \mem~190_q ;
wire \mem~222_q ;
wire \mem~158_q ;
wire \mem~336_combout ;
wire \mem~254_q ;
wire \mem~337_combout ;
wire \mem~94_q ;
wire \mem~62_q ;
wire \mem~30_q ;
wire \mem~338_combout ;
wire \mem~126_q ;
wire \mem~339_combout ;
wire \mem~340_combout ;
wire \internal_out_payload[30]~q ;
wire \mem~189_q ;
wire \mem~221_q ;
wire \mem~157_q ;
wire \mem~341_combout ;
wire \mem~253_q ;
wire \mem~342_combout ;
wire \mem~93_q ;
wire \mem~61_q ;
wire \mem~29_q ;
wire \mem~343_combout ;
wire \mem~125_q ;
wire \mem~344_combout ;
wire \mem~345_combout ;
wire \internal_out_payload[29]~q ;
wire \mem~188_q ;
wire \mem~220_q ;
wire \mem~156_q ;
wire \mem~346_combout ;
wire \mem~252_q ;
wire \mem~347_combout ;
wire \mem~92_q ;
wire \mem~60_q ;
wire \mem~28_q ;
wire \mem~348_combout ;
wire \mem~124_q ;
wire \mem~349_combout ;
wire \mem~350_combout ;
wire \internal_out_payload[28]~q ;
wire \mem~187_q ;
wire \mem~219_q ;
wire \mem~155_q ;
wire \mem~351_combout ;
wire \mem~251_q ;
wire \mem~352_combout ;
wire \mem~91_q ;
wire \mem~59_q ;
wire \mem~27_q ;
wire \mem~353_combout ;
wire \mem~123_q ;
wire \mem~354_combout ;
wire \mem~355_combout ;
wire \internal_out_payload[27]~q ;
wire \mem~186_q ;
wire \mem~218_q ;
wire \mem~154_q ;
wire \mem~356_combout ;
wire \mem~250_q ;
wire \mem~357_combout ;
wire \mem~90_q ;
wire \mem~58_q ;
wire \mem~26_q ;
wire \mem~358_combout ;
wire \mem~122_q ;
wire \mem~359_combout ;
wire \mem~360_combout ;
wire \internal_out_payload[26]~q ;
wire \mem~185_q ;
wire \mem~217_q ;
wire \mem~153_q ;
wire \mem~361_combout ;
wire \mem~249_q ;
wire \mem~362_combout ;
wire \mem~89_q ;
wire \mem~57_q ;
wire \mem~25_q ;
wire \mem~363_combout ;
wire \mem~121_q ;
wire \mem~364_combout ;
wire \mem~365_combout ;
wire \internal_out_payload[25]~q ;
wire \mem~170_q ;
wire \mem~202_q ;
wire \mem~138_q ;
wire \mem~366_combout ;
wire \mem~234_q ;
wire \mem~367_combout ;
wire \mem~74_q ;
wire \mem~42_q ;
wire \mem~10_q ;
wire \mem~368_combout ;
wire \mem~106_q ;
wire \mem~369_combout ;
wire \mem~370_combout ;
wire \internal_out_payload[10]~q ;
wire \mem~184_q ;
wire \mem~216_q ;
wire \mem~152_q ;
wire \mem~371_combout ;
wire \mem~248_q ;
wire \mem~372_combout ;
wire \mem~88_q ;
wire \mem~56_q ;
wire \mem~24_q ;
wire \mem~373_combout ;
wire \mem~120_q ;
wire \mem~374_combout ;
wire \mem~375_combout ;
wire \internal_out_payload[24]~q ;
wire \mem~169_q ;
wire \mem~201_q ;
wire \mem~137_q ;
wire \mem~376_combout ;
wire \mem~233_q ;
wire \mem~377_combout ;
wire \mem~73_q ;
wire \mem~41_q ;
wire \mem~9_q ;
wire \mem~378_combout ;
wire \mem~105_q ;
wire \mem~379_combout ;
wire \mem~380_combout ;
wire \internal_out_payload[9]~q ;
wire \mem~183_q ;
wire \mem~215_q ;
wire \mem~151_q ;
wire \mem~381_combout ;
wire \mem~247_q ;
wire \mem~382_combout ;
wire \mem~87_q ;
wire \mem~55_q ;
wire \mem~23_q ;
wire \mem~383_combout ;
wire \mem~119_q ;
wire \mem~384_combout ;
wire \mem~385_combout ;
wire \internal_out_payload[23]~q ;
wire \mem~168_q ;
wire \mem~200_q ;
wire \mem~136_q ;
wire \mem~386_combout ;
wire \mem~232_q ;
wire \mem~387_combout ;
wire \mem~72_q ;
wire \mem~40_q ;
wire \mem~8_q ;
wire \mem~388_combout ;
wire \mem~104_q ;
wire \mem~389_combout ;
wire \mem~390_combout ;
wire \internal_out_payload[8]~q ;
wire \mem~182_q ;
wire \mem~214_q ;
wire \mem~150_q ;
wire \mem~391_combout ;
wire \mem~246_q ;
wire \mem~392_combout ;
wire \mem~86_q ;
wire \mem~54_q ;
wire \mem~22_q ;
wire \mem~393_combout ;
wire \mem~118_q ;
wire \mem~394_combout ;
wire \mem~395_combout ;
wire \internal_out_payload[22]~q ;
wire \mem~167_q ;
wire \mem~199_q ;
wire \mem~135_q ;
wire \mem~396_combout ;
wire \mem~231_q ;
wire \mem~397_combout ;
wire \mem~71_q ;
wire \mem~39_q ;
wire \mem~7_q ;
wire \mem~398_combout ;
wire \mem~103_q ;
wire \mem~399_combout ;
wire \mem~400_combout ;
wire \internal_out_payload[7]~q ;
wire \mem~166_q ;
wire \mem~198_q ;
wire \mem~134_q ;
wire \mem~401_combout ;
wire \mem~230_q ;
wire \mem~402_combout ;
wire \mem~70_q ;
wire \mem~38_q ;
wire \mem~6_q ;
wire \mem~403_combout ;
wire \mem~102_q ;
wire \mem~404_combout ;
wire \mem~405_combout ;
wire \internal_out_payload[6]~q ;
wire \mem~180_q ;
wire \mem~212_q ;
wire \mem~148_q ;
wire \mem~406_combout ;
wire \mem~244_q ;
wire \mem~407_combout ;
wire \mem~84_q ;
wire \mem~52_q ;
wire \mem~20_q ;
wire \mem~408_combout ;
wire \mem~116_q ;
wire \mem~409_combout ;
wire \mem~410_combout ;
wire \internal_out_payload[20]~q ;
wire \mem~179_q ;
wire \mem~211_q ;
wire \mem~147_q ;
wire \mem~411_combout ;
wire \mem~243_q ;
wire \mem~412_combout ;
wire \mem~83_q ;
wire \mem~51_q ;
wire \mem~19_q ;
wire \mem~413_combout ;
wire \mem~115_q ;
wire \mem~414_combout ;
wire \mem~415_combout ;
wire \internal_out_payload[19]~q ;


dffeas out_valid(
	.clk(clk),
	.d(\internal_out_valid~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[0] (
	.clk(clk),
	.d(\internal_out_payload[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk),
	.d(\internal_out_payload[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk),
	.d(\internal_out_payload[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas \out_payload[3] (
	.clk(clk),
	.d(\internal_out_payload[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_3),
	.prn(vcc));
defparam \out_payload[3] .is_wysiwyg = "true";
defparam \out_payload[3] .power_up = "low";

dffeas \out_payload[4] (
	.clk(clk),
	.d(\internal_out_payload[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_4),
	.prn(vcc));
defparam \out_payload[4] .is_wysiwyg = "true";
defparam \out_payload[4] .power_up = "low";

dffeas \out_payload[11] (
	.clk(clk),
	.d(\internal_out_payload[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_11),
	.prn(vcc));
defparam \out_payload[11] .is_wysiwyg = "true";
defparam \out_payload[11] .power_up = "low";

dffeas \out_payload[13] (
	.clk(clk),
	.d(\internal_out_payload[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_13),
	.prn(vcc));
defparam \out_payload[13] .is_wysiwyg = "true";
defparam \out_payload[13] .power_up = "low";

dffeas \out_payload[16] (
	.clk(clk),
	.d(\internal_out_payload[16]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_16),
	.prn(vcc));
defparam \out_payload[16] .is_wysiwyg = "true";
defparam \out_payload[16] .power_up = "low";

dffeas \out_payload[12] (
	.clk(clk),
	.d(\internal_out_payload[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[5] (
	.clk(clk),
	.d(\internal_out_payload[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[14] (
	.clk(clk),
	.d(\internal_out_payload[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_14),
	.prn(vcc));
defparam \out_payload[14] .is_wysiwyg = "true";
defparam \out_payload[14] .power_up = "low";

dffeas \out_payload[15] (
	.clk(clk),
	.d(\internal_out_payload[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_15),
	.prn(vcc));
defparam \out_payload[15] .is_wysiwyg = "true";
defparam \out_payload[15] .power_up = "low";

dffeas \out_payload[21] (
	.clk(clk),
	.d(\internal_out_payload[21]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_21),
	.prn(vcc));
defparam \out_payload[21] .is_wysiwyg = "true";
defparam \out_payload[21] .power_up = "low";

dffeas \out_payload[18] (
	.clk(clk),
	.d(\internal_out_payload[18]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_18),
	.prn(vcc));
defparam \out_payload[18] .is_wysiwyg = "true";
defparam \out_payload[18] .power_up = "low";

dffeas \out_payload[17] (
	.clk(clk),
	.d(\internal_out_payload[17]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_17),
	.prn(vcc));
defparam \out_payload[17] .is_wysiwyg = "true";
defparam \out_payload[17] .power_up = "low";

dffeas \out_payload[31] (
	.clk(clk),
	.d(\internal_out_payload[31]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_31),
	.prn(vcc));
defparam \out_payload[31] .is_wysiwyg = "true";
defparam \out_payload[31] .power_up = "low";

dffeas \out_payload[30] (
	.clk(clk),
	.d(\internal_out_payload[30]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_30),
	.prn(vcc));
defparam \out_payload[30] .is_wysiwyg = "true";
defparam \out_payload[30] .power_up = "low";

dffeas \out_payload[29] (
	.clk(clk),
	.d(\internal_out_payload[29]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_29),
	.prn(vcc));
defparam \out_payload[29] .is_wysiwyg = "true";
defparam \out_payload[29] .power_up = "low";

dffeas \out_payload[28] (
	.clk(clk),
	.d(\internal_out_payload[28]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_28),
	.prn(vcc));
defparam \out_payload[28] .is_wysiwyg = "true";
defparam \out_payload[28] .power_up = "low";

dffeas \out_payload[27] (
	.clk(clk),
	.d(\internal_out_payload[27]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_27),
	.prn(vcc));
defparam \out_payload[27] .is_wysiwyg = "true";
defparam \out_payload[27] .power_up = "low";

dffeas \out_payload[26] (
	.clk(clk),
	.d(\internal_out_payload[26]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_26),
	.prn(vcc));
defparam \out_payload[26] .is_wysiwyg = "true";
defparam \out_payload[26] .power_up = "low";

dffeas \out_payload[25] (
	.clk(clk),
	.d(\internal_out_payload[25]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_25),
	.prn(vcc));
defparam \out_payload[25] .is_wysiwyg = "true";
defparam \out_payload[25] .power_up = "low";

dffeas \out_payload[10] (
	.clk(clk),
	.d(\internal_out_payload[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_10),
	.prn(vcc));
defparam \out_payload[10] .is_wysiwyg = "true";
defparam \out_payload[10] .power_up = "low";

dffeas \out_payload[24] (
	.clk(clk),
	.d(\internal_out_payload[24]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_24),
	.prn(vcc));
defparam \out_payload[24] .is_wysiwyg = "true";
defparam \out_payload[24] .power_up = "low";

dffeas \out_payload[9] (
	.clk(clk),
	.d(\internal_out_payload[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_9),
	.prn(vcc));
defparam \out_payload[9] .is_wysiwyg = "true";
defparam \out_payload[9] .power_up = "low";

dffeas \out_payload[23] (
	.clk(clk),
	.d(\internal_out_payload[23]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_23),
	.prn(vcc));
defparam \out_payload[23] .is_wysiwyg = "true";
defparam \out_payload[23] .power_up = "low";

dffeas \out_payload[8] (
	.clk(clk),
	.d(\internal_out_payload[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

dffeas \out_payload[22] (
	.clk(clk),
	.d(\internal_out_payload[22]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_22),
	.prn(vcc));
defparam \out_payload[22] .is_wysiwyg = "true";
defparam \out_payload[22] .power_up = "low";

dffeas \out_payload[7] (
	.clk(clk),
	.d(\internal_out_payload[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[6] (
	.clk(clk),
	.d(\internal_out_payload[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

dffeas \out_payload[20] (
	.clk(clk),
	.d(\internal_out_payload[20]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_20),
	.prn(vcc));
defparam \out_payload[20] .is_wysiwyg = "true";
defparam \out_payload[20] .power_up = "low";

dffeas \out_payload[19] (
	.clk(clk),
	.d(\internal_out_payload[19]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~0_combout ),
	.q(out_payload_19),
	.prn(vcc));
defparam \out_payload[19] .is_wysiwyg = "true";
defparam \out_payload[19] .power_up = "low";

cycloneive_lcell_comb \internal_out_ready~0 (
	.dataa(mem_used_0),
	.datab(mem_107_0),
	.datac(WideOr0),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_ready~0_combout ),
	.cout());
defparam \internal_out_ready~0 .lut_mask = 16'h7FFF;
defparam \internal_out_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[0]~1 (
	.dataa(gnd),
	.datab(\rd_ptr[0]~q ),
	.datac(\internal_out_valid~q ),
	.datad(\internal_out_ready~0_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[0]~1_combout ),
	.cout());
defparam \mem_rd_ptr[0]~1 .lut_mask = 16'hC33C;
defparam \mem_rd_ptr[0]~1 .sum_lutc_input = "datac";

dffeas \rd_ptr[0] (
	.clk(clk),
	.d(\mem_rd_ptr[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[0]~q ),
	.prn(vcc));
defparam \rd_ptr[0] .is_wysiwyg = "true";
defparam \rd_ptr[0] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[1]~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\internal_out_valid~q ),
	.datac(\internal_out_ready~0_combout ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[1]~0_combout ),
	.cout());
defparam \mem_rd_ptr[1]~0 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[1]~0 .sum_lutc_input = "datac";

dffeas \rd_ptr[1] (
	.clk(clk),
	.d(\mem_rd_ptr[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[1]~q ),
	.prn(vcc));
defparam \rd_ptr[1] .is_wysiwyg = "true";
defparam \rd_ptr[1] .power_up = "low";

cycloneive_lcell_comb \wr_ptr[0]~0 (
	.dataa(\wr_ptr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_ptr[0]~0_combout ),
	.cout());
defparam \wr_ptr[0]~0 .lut_mask = 16'h5555;
defparam \wr_ptr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\next_full~0_combout ),
	.cout());
defparam \next_full~0 .lut_mask = 16'h6996;
defparam \next_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(\internal_out_valid~q ),
	.datab(\internal_out_ready~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hEEEE;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[2]~2 (
	.dataa(\rd_ptr[2]~q ),
	.datab(\read~0_combout ),
	.datac(\rd_ptr[1]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[2]~2_combout ),
	.cout());
defparam \mem_rd_ptr[2]~2 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[2]~2 .sum_lutc_input = "datac";

dffeas \rd_ptr[2] (
	.clk(clk),
	.d(\mem_rd_ptr[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[2]~q ),
	.prn(vcc));
defparam \rd_ptr[2] .is_wysiwyg = "true";
defparam \rd_ptr[2] .power_up = "low";

dffeas \wr_ptr[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_ptr[2] .is_wysiwyg = "true";
defparam \wr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'hC33C;
defparam \Add0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~1 (
	.dataa(za_valid),
	.datab(\next_full~0_combout ),
	.datac(\rd_ptr[2]~q ),
	.datad(\Add0~1_combout ),
	.cin(gnd),
	.combout(\next_full~1_combout ),
	.cout());
defparam \next_full~1 .lut_mask = 16'hEFFE;
defparam \next_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~2 (
	.dataa(\full~q ),
	.datab(\next_full~1_combout ),
	.datac(\internal_out_valid~q ),
	.datad(\internal_out_ready~0_combout ),
	.cin(gnd),
	.combout(\next_full~2_combout ),
	.cout());
defparam \next_full~2 .lut_mask = 16'hEFFF;
defparam \next_full~2 .sum_lutc_input = "datac";

dffeas full(
	.clk(clk),
	.d(\next_full~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\full~q ),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

cycloneive_lcell_comb write(
	.dataa(za_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(\full~q ),
	.cin(gnd),
	.combout(\write~combout ),
	.cout());
defparam write.lut_mask = 16'hAAFF;
defparam write.sum_lutc_input = "datac";

dffeas \wr_ptr[0] (
	.clk(clk),
	.d(\wr_ptr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_ptr[0] .is_wysiwyg = "true";
defparam \wr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \wr_ptr[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_ptr[1] .is_wysiwyg = "true";
defparam \wr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \internal_out_valid~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\internal_out_valid~0_combout ),
	.cout());
defparam \internal_out_valid~0 .lut_mask = 16'h6996;
defparam \internal_out_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\rd_ptr[0]~q ),
	.datac(\wr_ptr[2]~q ),
	.datad(\rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_valid~1 (
	.dataa(\internal_out_valid~q ),
	.datab(\internal_out_ready~0_combout ),
	.datac(\internal_out_valid~0_combout ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~1_combout ),
	.cout());
defparam \internal_out_valid~1 .lut_mask = 16'hFEFF;
defparam \internal_out_valid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_empty~0 (
	.dataa(\read~0_combout ),
	.datab(\internal_out_valid~1_combout ),
	.datac(\empty~q ),
	.datad(\write~combout ),
	.cin(gnd),
	.combout(\next_empty~0_combout ),
	.cout());
defparam \next_empty~0 .lut_mask = 16'hFFF7;
defparam \next_empty~0 .sum_lutc_input = "datac";

dffeas empty(
	.clk(clk),
	.d(\next_empty~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

cycloneive_lcell_comb \internal_out_valid~2 (
	.dataa(\internal_out_valid~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\empty~q ),
	.cin(gnd),
	.combout(\internal_out_valid~2_combout ),
	.cout());
defparam \internal_out_valid~2 .lut_mask = 16'hFF55;
defparam \internal_out_valid~2 .sum_lutc_input = "datac";

dffeas internal_out_valid(
	.clk(clk),
	.d(\internal_out_valid~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_valid~q ),
	.prn(vcc));
defparam internal_out_valid.is_wysiwyg = "true";
defparam internal_out_valid.power_up = "low";

cycloneive_lcell_comb \mem~416 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~416_combout ),
	.cout());
defparam \mem~416 .lut_mask = 16'hFEFF;
defparam \mem~416 .sum_lutc_input = "datac";

dffeas \mem~160 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~160_q ),
	.prn(vcc));
defparam \mem~160 .is_wysiwyg = "true";
defparam \mem~160 .power_up = "low";

cycloneive_lcell_comb \mem~417 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem~417_combout ),
	.cout());
defparam \mem~417 .lut_mask = 16'hFEFF;
defparam \mem~417 .sum_lutc_input = "datac";

dffeas \mem~192 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~192_q ),
	.prn(vcc));
defparam \mem~192 .is_wysiwyg = "true";
defparam \mem~192 .power_up = "low";

cycloneive_lcell_comb \mem~418 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~418_combout ),
	.cout());
defparam \mem~418 .lut_mask = 16'hEFFF;
defparam \mem~418 .sum_lutc_input = "datac";

dffeas \mem~128 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~128_q ),
	.prn(vcc));
defparam \mem~128 .is_wysiwyg = "true";
defparam \mem~128 .power_up = "low";

cycloneive_lcell_comb \mem~256 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~192_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~128_q ),
	.cin(gnd),
	.combout(\mem~256_combout ),
	.cout());
defparam \mem~256 .lut_mask = 16'hFFDE;
defparam \mem~256 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~419 (
	.dataa(\wr_ptr[2]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\write~combout ),
	.cin(gnd),
	.combout(\mem~419_combout ),
	.cout());
defparam \mem~419 .lut_mask = 16'hFFFE;
defparam \mem~419 .sum_lutc_input = "datac";

dffeas \mem~224 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~224_q ),
	.prn(vcc));
defparam \mem~224 .is_wysiwyg = "true";
defparam \mem~224 .power_up = "low";

cycloneive_lcell_comb \mem~257 (
	.dataa(\mem~160_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~256_combout ),
	.datad(\mem~224_q ),
	.cin(gnd),
	.combout(\mem~257_combout ),
	.cout());
defparam \mem~257 .lut_mask = 16'hFFBE;
defparam \mem~257 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~420 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem~420_combout ),
	.cout());
defparam \mem~420 .lut_mask = 16'hEFFF;
defparam \mem~420 .sum_lutc_input = "datac";

dffeas \mem~64 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~64_q ),
	.prn(vcc));
defparam \mem~64 .is_wysiwyg = "true";
defparam \mem~64 .power_up = "low";

cycloneive_lcell_comb \mem~421 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\write~combout ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~421_combout ),
	.cout());
defparam \mem~421 .lut_mask = 16'hEFFF;
defparam \mem~421 .sum_lutc_input = "datac";

dffeas \mem~32 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~32_q ),
	.prn(vcc));
defparam \mem~32 .is_wysiwyg = "true";
defparam \mem~32 .power_up = "low";

cycloneive_lcell_comb \mem~422 (
	.dataa(\write~combout ),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem~422_combout ),
	.cout());
defparam \mem~422 .lut_mask = 16'hBFFF;
defparam \mem~422 .sum_lutc_input = "datac";

dffeas \mem~0 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~0_q ),
	.prn(vcc));
defparam \mem~0 .is_wysiwyg = "true";
defparam \mem~0 .power_up = "low";

cycloneive_lcell_comb \mem~258 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~32_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~0_q ),
	.cin(gnd),
	.combout(\mem~258_combout ),
	.cout());
defparam \mem~258 .lut_mask = 16'hFFDE;
defparam \mem~258 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~423 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\write~combout ),
	.datad(\wr_ptr[2]~q ),
	.cin(gnd),
	.combout(\mem~423_combout ),
	.cout());
defparam \mem~423 .lut_mask = 16'hFEFF;
defparam \mem~423 .sum_lutc_input = "datac";

dffeas \mem~96 (
	.clk(clk),
	.d(za_data_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~96_q ),
	.prn(vcc));
defparam \mem~96 .is_wysiwyg = "true";
defparam \mem~96 .power_up = "low";

cycloneive_lcell_comb \mem~259 (
	.dataa(\mem~64_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~258_combout ),
	.datad(\mem~96_q ),
	.cin(gnd),
	.combout(\mem~259_combout ),
	.cout());
defparam \mem~259 .lut_mask = 16'hFFBE;
defparam \mem~259 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~260 (
	.dataa(\mem~257_combout ),
	.datab(\mem~259_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~260_combout ),
	.cout());
defparam \mem~260 .lut_mask = 16'hAACC;
defparam \mem~260 .sum_lutc_input = "datac";

dffeas \internal_out_payload[0] (
	.clk(clk),
	.d(\mem~260_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[0]~q ),
	.prn(vcc));
defparam \internal_out_payload[0] .is_wysiwyg = "true";
defparam \internal_out_payload[0] .power_up = "low";

dffeas \mem~161 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~161_q ),
	.prn(vcc));
defparam \mem~161 .is_wysiwyg = "true";
defparam \mem~161 .power_up = "low";

dffeas \mem~193 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~193_q ),
	.prn(vcc));
defparam \mem~193 .is_wysiwyg = "true";
defparam \mem~193 .power_up = "low";

dffeas \mem~129 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~129_q ),
	.prn(vcc));
defparam \mem~129 .is_wysiwyg = "true";
defparam \mem~129 .power_up = "low";

cycloneive_lcell_comb \mem~261 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~193_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~129_q ),
	.cin(gnd),
	.combout(\mem~261_combout ),
	.cout());
defparam \mem~261 .lut_mask = 16'hFFDE;
defparam \mem~261 .sum_lutc_input = "datac";

dffeas \mem~225 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~225_q ),
	.prn(vcc));
defparam \mem~225 .is_wysiwyg = "true";
defparam \mem~225 .power_up = "low";

cycloneive_lcell_comb \mem~262 (
	.dataa(\mem~161_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~261_combout ),
	.datad(\mem~225_q ),
	.cin(gnd),
	.combout(\mem~262_combout ),
	.cout());
defparam \mem~262 .lut_mask = 16'hFFBE;
defparam \mem~262 .sum_lutc_input = "datac";

dffeas \mem~65 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~65_q ),
	.prn(vcc));
defparam \mem~65 .is_wysiwyg = "true";
defparam \mem~65 .power_up = "low";

dffeas \mem~33 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~33_q ),
	.prn(vcc));
defparam \mem~33 .is_wysiwyg = "true";
defparam \mem~33 .power_up = "low";

dffeas \mem~1 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~1_q ),
	.prn(vcc));
defparam \mem~1 .is_wysiwyg = "true";
defparam \mem~1 .power_up = "low";

cycloneive_lcell_comb \mem~263 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~33_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~1_q ),
	.cin(gnd),
	.combout(\mem~263_combout ),
	.cout());
defparam \mem~263 .lut_mask = 16'hFFDE;
defparam \mem~263 .sum_lutc_input = "datac";

dffeas \mem~97 (
	.clk(clk),
	.d(za_data_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~97_q ),
	.prn(vcc));
defparam \mem~97 .is_wysiwyg = "true";
defparam \mem~97 .power_up = "low";

cycloneive_lcell_comb \mem~264 (
	.dataa(\mem~65_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~263_combout ),
	.datad(\mem~97_q ),
	.cin(gnd),
	.combout(\mem~264_combout ),
	.cout());
defparam \mem~264 .lut_mask = 16'hFFBE;
defparam \mem~264 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~265 (
	.dataa(\mem~262_combout ),
	.datab(\mem~264_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~265_combout ),
	.cout());
defparam \mem~265 .lut_mask = 16'hAACC;
defparam \mem~265 .sum_lutc_input = "datac";

dffeas \internal_out_payload[1] (
	.clk(clk),
	.d(\mem~265_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[1]~q ),
	.prn(vcc));
defparam \internal_out_payload[1] .is_wysiwyg = "true";
defparam \internal_out_payload[1] .power_up = "low";

dffeas \mem~162 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~162_q ),
	.prn(vcc));
defparam \mem~162 .is_wysiwyg = "true";
defparam \mem~162 .power_up = "low";

dffeas \mem~194 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~194_q ),
	.prn(vcc));
defparam \mem~194 .is_wysiwyg = "true";
defparam \mem~194 .power_up = "low";

dffeas \mem~130 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~130_q ),
	.prn(vcc));
defparam \mem~130 .is_wysiwyg = "true";
defparam \mem~130 .power_up = "low";

cycloneive_lcell_comb \mem~266 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~194_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~130_q ),
	.cin(gnd),
	.combout(\mem~266_combout ),
	.cout());
defparam \mem~266 .lut_mask = 16'hFFDE;
defparam \mem~266 .sum_lutc_input = "datac";

dffeas \mem~226 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~226_q ),
	.prn(vcc));
defparam \mem~226 .is_wysiwyg = "true";
defparam \mem~226 .power_up = "low";

cycloneive_lcell_comb \mem~267 (
	.dataa(\mem~162_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~266_combout ),
	.datad(\mem~226_q ),
	.cin(gnd),
	.combout(\mem~267_combout ),
	.cout());
defparam \mem~267 .lut_mask = 16'hFFBE;
defparam \mem~267 .sum_lutc_input = "datac";

dffeas \mem~66 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~66_q ),
	.prn(vcc));
defparam \mem~66 .is_wysiwyg = "true";
defparam \mem~66 .power_up = "low";

dffeas \mem~34 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~34_q ),
	.prn(vcc));
defparam \mem~34 .is_wysiwyg = "true";
defparam \mem~34 .power_up = "low";

dffeas \mem~2 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~2_q ),
	.prn(vcc));
defparam \mem~2 .is_wysiwyg = "true";
defparam \mem~2 .power_up = "low";

cycloneive_lcell_comb \mem~268 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~34_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~2_q ),
	.cin(gnd),
	.combout(\mem~268_combout ),
	.cout());
defparam \mem~268 .lut_mask = 16'hFFDE;
defparam \mem~268 .sum_lutc_input = "datac";

dffeas \mem~98 (
	.clk(clk),
	.d(za_data_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~98_q ),
	.prn(vcc));
defparam \mem~98 .is_wysiwyg = "true";
defparam \mem~98 .power_up = "low";

cycloneive_lcell_comb \mem~269 (
	.dataa(\mem~66_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~268_combout ),
	.datad(\mem~98_q ),
	.cin(gnd),
	.combout(\mem~269_combout ),
	.cout());
defparam \mem~269 .lut_mask = 16'hFFBE;
defparam \mem~269 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~270 (
	.dataa(\mem~267_combout ),
	.datab(\mem~269_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~270_combout ),
	.cout());
defparam \mem~270 .lut_mask = 16'hAACC;
defparam \mem~270 .sum_lutc_input = "datac";

dffeas \internal_out_payload[2] (
	.clk(clk),
	.d(\mem~270_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[2]~q ),
	.prn(vcc));
defparam \internal_out_payload[2] .is_wysiwyg = "true";
defparam \internal_out_payload[2] .power_up = "low";

dffeas \mem~163 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~163_q ),
	.prn(vcc));
defparam \mem~163 .is_wysiwyg = "true";
defparam \mem~163 .power_up = "low";

dffeas \mem~195 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~195_q ),
	.prn(vcc));
defparam \mem~195 .is_wysiwyg = "true";
defparam \mem~195 .power_up = "low";

dffeas \mem~131 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~131_q ),
	.prn(vcc));
defparam \mem~131 .is_wysiwyg = "true";
defparam \mem~131 .power_up = "low";

cycloneive_lcell_comb \mem~271 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~195_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~131_q ),
	.cin(gnd),
	.combout(\mem~271_combout ),
	.cout());
defparam \mem~271 .lut_mask = 16'hFFDE;
defparam \mem~271 .sum_lutc_input = "datac";

dffeas \mem~227 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~227_q ),
	.prn(vcc));
defparam \mem~227 .is_wysiwyg = "true";
defparam \mem~227 .power_up = "low";

cycloneive_lcell_comb \mem~272 (
	.dataa(\mem~163_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~271_combout ),
	.datad(\mem~227_q ),
	.cin(gnd),
	.combout(\mem~272_combout ),
	.cout());
defparam \mem~272 .lut_mask = 16'hFFBE;
defparam \mem~272 .sum_lutc_input = "datac";

dffeas \mem~67 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~67_q ),
	.prn(vcc));
defparam \mem~67 .is_wysiwyg = "true";
defparam \mem~67 .power_up = "low";

dffeas \mem~35 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~35_q ),
	.prn(vcc));
defparam \mem~35 .is_wysiwyg = "true";
defparam \mem~35 .power_up = "low";

dffeas \mem~3 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~3_q ),
	.prn(vcc));
defparam \mem~3 .is_wysiwyg = "true";
defparam \mem~3 .power_up = "low";

cycloneive_lcell_comb \mem~273 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~35_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~3_q ),
	.cin(gnd),
	.combout(\mem~273_combout ),
	.cout());
defparam \mem~273 .lut_mask = 16'hFFDE;
defparam \mem~273 .sum_lutc_input = "datac";

dffeas \mem~99 (
	.clk(clk),
	.d(za_data_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~99_q ),
	.prn(vcc));
defparam \mem~99 .is_wysiwyg = "true";
defparam \mem~99 .power_up = "low";

cycloneive_lcell_comb \mem~274 (
	.dataa(\mem~67_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~273_combout ),
	.datad(\mem~99_q ),
	.cin(gnd),
	.combout(\mem~274_combout ),
	.cout());
defparam \mem~274 .lut_mask = 16'hFFBE;
defparam \mem~274 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~275 (
	.dataa(\mem~272_combout ),
	.datab(\mem~274_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~275_combout ),
	.cout());
defparam \mem~275 .lut_mask = 16'hAACC;
defparam \mem~275 .sum_lutc_input = "datac";

dffeas \internal_out_payload[3] (
	.clk(clk),
	.d(\mem~275_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[3]~q ),
	.prn(vcc));
defparam \internal_out_payload[3] .is_wysiwyg = "true";
defparam \internal_out_payload[3] .power_up = "low";

dffeas \mem~164 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~164_q ),
	.prn(vcc));
defparam \mem~164 .is_wysiwyg = "true";
defparam \mem~164 .power_up = "low";

dffeas \mem~196 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~196_q ),
	.prn(vcc));
defparam \mem~196 .is_wysiwyg = "true";
defparam \mem~196 .power_up = "low";

dffeas \mem~132 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~132_q ),
	.prn(vcc));
defparam \mem~132 .is_wysiwyg = "true";
defparam \mem~132 .power_up = "low";

cycloneive_lcell_comb \mem~276 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~196_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~132_q ),
	.cin(gnd),
	.combout(\mem~276_combout ),
	.cout());
defparam \mem~276 .lut_mask = 16'hFFDE;
defparam \mem~276 .sum_lutc_input = "datac";

dffeas \mem~228 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~228_q ),
	.prn(vcc));
defparam \mem~228 .is_wysiwyg = "true";
defparam \mem~228 .power_up = "low";

cycloneive_lcell_comb \mem~277 (
	.dataa(\mem~164_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~276_combout ),
	.datad(\mem~228_q ),
	.cin(gnd),
	.combout(\mem~277_combout ),
	.cout());
defparam \mem~277 .lut_mask = 16'hFFBE;
defparam \mem~277 .sum_lutc_input = "datac";

dffeas \mem~68 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~68_q ),
	.prn(vcc));
defparam \mem~68 .is_wysiwyg = "true";
defparam \mem~68 .power_up = "low";

dffeas \mem~36 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~36_q ),
	.prn(vcc));
defparam \mem~36 .is_wysiwyg = "true";
defparam \mem~36 .power_up = "low";

dffeas \mem~4 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~4_q ),
	.prn(vcc));
defparam \mem~4 .is_wysiwyg = "true";
defparam \mem~4 .power_up = "low";

cycloneive_lcell_comb \mem~278 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~36_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~4_q ),
	.cin(gnd),
	.combout(\mem~278_combout ),
	.cout());
defparam \mem~278 .lut_mask = 16'hFFDE;
defparam \mem~278 .sum_lutc_input = "datac";

dffeas \mem~100 (
	.clk(clk),
	.d(za_data_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~100_q ),
	.prn(vcc));
defparam \mem~100 .is_wysiwyg = "true";
defparam \mem~100 .power_up = "low";

cycloneive_lcell_comb \mem~279 (
	.dataa(\mem~68_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~278_combout ),
	.datad(\mem~100_q ),
	.cin(gnd),
	.combout(\mem~279_combout ),
	.cout());
defparam \mem~279 .lut_mask = 16'hFFBE;
defparam \mem~279 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~280 (
	.dataa(\mem~277_combout ),
	.datab(\mem~279_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~280_combout ),
	.cout());
defparam \mem~280 .lut_mask = 16'hAACC;
defparam \mem~280 .sum_lutc_input = "datac";

dffeas \internal_out_payload[4] (
	.clk(clk),
	.d(\mem~280_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[4]~q ),
	.prn(vcc));
defparam \internal_out_payload[4] .is_wysiwyg = "true";
defparam \internal_out_payload[4] .power_up = "low";

dffeas \mem~171 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~171_q ),
	.prn(vcc));
defparam \mem~171 .is_wysiwyg = "true";
defparam \mem~171 .power_up = "low";

dffeas \mem~203 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~203_q ),
	.prn(vcc));
defparam \mem~203 .is_wysiwyg = "true";
defparam \mem~203 .power_up = "low";

dffeas \mem~139 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~139_q ),
	.prn(vcc));
defparam \mem~139 .is_wysiwyg = "true";
defparam \mem~139 .power_up = "low";

cycloneive_lcell_comb \mem~281 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~203_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~139_q ),
	.cin(gnd),
	.combout(\mem~281_combout ),
	.cout());
defparam \mem~281 .lut_mask = 16'hFFDE;
defparam \mem~281 .sum_lutc_input = "datac";

dffeas \mem~235 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~235_q ),
	.prn(vcc));
defparam \mem~235 .is_wysiwyg = "true";
defparam \mem~235 .power_up = "low";

cycloneive_lcell_comb \mem~282 (
	.dataa(\mem~171_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~281_combout ),
	.datad(\mem~235_q ),
	.cin(gnd),
	.combout(\mem~282_combout ),
	.cout());
defparam \mem~282 .lut_mask = 16'hFFBE;
defparam \mem~282 .sum_lutc_input = "datac";

dffeas \mem~75 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~75_q ),
	.prn(vcc));
defparam \mem~75 .is_wysiwyg = "true";
defparam \mem~75 .power_up = "low";

dffeas \mem~43 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~43_q ),
	.prn(vcc));
defparam \mem~43 .is_wysiwyg = "true";
defparam \mem~43 .power_up = "low";

dffeas \mem~11 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~11_q ),
	.prn(vcc));
defparam \mem~11 .is_wysiwyg = "true";
defparam \mem~11 .power_up = "low";

cycloneive_lcell_comb \mem~283 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~43_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~11_q ),
	.cin(gnd),
	.combout(\mem~283_combout ),
	.cout());
defparam \mem~283 .lut_mask = 16'hFFDE;
defparam \mem~283 .sum_lutc_input = "datac";

dffeas \mem~107 (
	.clk(clk),
	.d(za_data_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~107_q ),
	.prn(vcc));
defparam \mem~107 .is_wysiwyg = "true";
defparam \mem~107 .power_up = "low";

cycloneive_lcell_comb \mem~284 (
	.dataa(\mem~75_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~283_combout ),
	.datad(\mem~107_q ),
	.cin(gnd),
	.combout(\mem~284_combout ),
	.cout());
defparam \mem~284 .lut_mask = 16'hFFBE;
defparam \mem~284 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~285 (
	.dataa(\mem~282_combout ),
	.datab(\mem~284_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~285_combout ),
	.cout());
defparam \mem~285 .lut_mask = 16'hAACC;
defparam \mem~285 .sum_lutc_input = "datac";

dffeas \internal_out_payload[11] (
	.clk(clk),
	.d(\mem~285_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[11]~q ),
	.prn(vcc));
defparam \internal_out_payload[11] .is_wysiwyg = "true";
defparam \internal_out_payload[11] .power_up = "low";

dffeas \mem~173 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~173_q ),
	.prn(vcc));
defparam \mem~173 .is_wysiwyg = "true";
defparam \mem~173 .power_up = "low";

dffeas \mem~205 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~205_q ),
	.prn(vcc));
defparam \mem~205 .is_wysiwyg = "true";
defparam \mem~205 .power_up = "low";

dffeas \mem~141 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~141_q ),
	.prn(vcc));
defparam \mem~141 .is_wysiwyg = "true";
defparam \mem~141 .power_up = "low";

cycloneive_lcell_comb \mem~286 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~205_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~141_q ),
	.cin(gnd),
	.combout(\mem~286_combout ),
	.cout());
defparam \mem~286 .lut_mask = 16'hFFDE;
defparam \mem~286 .sum_lutc_input = "datac";

dffeas \mem~237 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~237_q ),
	.prn(vcc));
defparam \mem~237 .is_wysiwyg = "true";
defparam \mem~237 .power_up = "low";

cycloneive_lcell_comb \mem~287 (
	.dataa(\mem~173_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~286_combout ),
	.datad(\mem~237_q ),
	.cin(gnd),
	.combout(\mem~287_combout ),
	.cout());
defparam \mem~287 .lut_mask = 16'hFFBE;
defparam \mem~287 .sum_lutc_input = "datac";

dffeas \mem~77 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~77_q ),
	.prn(vcc));
defparam \mem~77 .is_wysiwyg = "true";
defparam \mem~77 .power_up = "low";

dffeas \mem~45 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~45_q ),
	.prn(vcc));
defparam \mem~45 .is_wysiwyg = "true";
defparam \mem~45 .power_up = "low";

dffeas \mem~13 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~13_q ),
	.prn(vcc));
defparam \mem~13 .is_wysiwyg = "true";
defparam \mem~13 .power_up = "low";

cycloneive_lcell_comb \mem~288 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~45_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~13_q ),
	.cin(gnd),
	.combout(\mem~288_combout ),
	.cout());
defparam \mem~288 .lut_mask = 16'hFFDE;
defparam \mem~288 .sum_lutc_input = "datac";

dffeas \mem~109 (
	.clk(clk),
	.d(za_data_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~109_q ),
	.prn(vcc));
defparam \mem~109 .is_wysiwyg = "true";
defparam \mem~109 .power_up = "low";

cycloneive_lcell_comb \mem~289 (
	.dataa(\mem~77_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~288_combout ),
	.datad(\mem~109_q ),
	.cin(gnd),
	.combout(\mem~289_combout ),
	.cout());
defparam \mem~289 .lut_mask = 16'hFFBE;
defparam \mem~289 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~290 (
	.dataa(\mem~287_combout ),
	.datab(\mem~289_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~290_combout ),
	.cout());
defparam \mem~290 .lut_mask = 16'hAACC;
defparam \mem~290 .sum_lutc_input = "datac";

dffeas \internal_out_payload[13] (
	.clk(clk),
	.d(\mem~290_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[13]~q ),
	.prn(vcc));
defparam \internal_out_payload[13] .is_wysiwyg = "true";
defparam \internal_out_payload[13] .power_up = "low";

dffeas \mem~176 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~176_q ),
	.prn(vcc));
defparam \mem~176 .is_wysiwyg = "true";
defparam \mem~176 .power_up = "low";

dffeas \mem~208 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~208_q ),
	.prn(vcc));
defparam \mem~208 .is_wysiwyg = "true";
defparam \mem~208 .power_up = "low";

dffeas \mem~144 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~144_q ),
	.prn(vcc));
defparam \mem~144 .is_wysiwyg = "true";
defparam \mem~144 .power_up = "low";

cycloneive_lcell_comb \mem~291 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~208_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~144_q ),
	.cin(gnd),
	.combout(\mem~291_combout ),
	.cout());
defparam \mem~291 .lut_mask = 16'hFFDE;
defparam \mem~291 .sum_lutc_input = "datac";

dffeas \mem~240 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~240_q ),
	.prn(vcc));
defparam \mem~240 .is_wysiwyg = "true";
defparam \mem~240 .power_up = "low";

cycloneive_lcell_comb \mem~292 (
	.dataa(\mem~176_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~291_combout ),
	.datad(\mem~240_q ),
	.cin(gnd),
	.combout(\mem~292_combout ),
	.cout());
defparam \mem~292 .lut_mask = 16'hFFBE;
defparam \mem~292 .sum_lutc_input = "datac";

dffeas \mem~80 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~80_q ),
	.prn(vcc));
defparam \mem~80 .is_wysiwyg = "true";
defparam \mem~80 .power_up = "low";

dffeas \mem~48 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~48_q ),
	.prn(vcc));
defparam \mem~48 .is_wysiwyg = "true";
defparam \mem~48 .power_up = "low";

dffeas \mem~16 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~16_q ),
	.prn(vcc));
defparam \mem~16 .is_wysiwyg = "true";
defparam \mem~16 .power_up = "low";

cycloneive_lcell_comb \mem~293 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~48_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~16_q ),
	.cin(gnd),
	.combout(\mem~293_combout ),
	.cout());
defparam \mem~293 .lut_mask = 16'hFFDE;
defparam \mem~293 .sum_lutc_input = "datac";

dffeas \mem~112 (
	.clk(clk),
	.d(za_data_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~112_q ),
	.prn(vcc));
defparam \mem~112 .is_wysiwyg = "true";
defparam \mem~112 .power_up = "low";

cycloneive_lcell_comb \mem~294 (
	.dataa(\mem~80_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~293_combout ),
	.datad(\mem~112_q ),
	.cin(gnd),
	.combout(\mem~294_combout ),
	.cout());
defparam \mem~294 .lut_mask = 16'hFFBE;
defparam \mem~294 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~295 (
	.dataa(\mem~292_combout ),
	.datab(\mem~294_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~295_combout ),
	.cout());
defparam \mem~295 .lut_mask = 16'hAACC;
defparam \mem~295 .sum_lutc_input = "datac";

dffeas \internal_out_payload[16] (
	.clk(clk),
	.d(\mem~295_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[16]~q ),
	.prn(vcc));
defparam \internal_out_payload[16] .is_wysiwyg = "true";
defparam \internal_out_payload[16] .power_up = "low";

dffeas \mem~172 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~172_q ),
	.prn(vcc));
defparam \mem~172 .is_wysiwyg = "true";
defparam \mem~172 .power_up = "low";

dffeas \mem~204 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~204_q ),
	.prn(vcc));
defparam \mem~204 .is_wysiwyg = "true";
defparam \mem~204 .power_up = "low";

dffeas \mem~140 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~140_q ),
	.prn(vcc));
defparam \mem~140 .is_wysiwyg = "true";
defparam \mem~140 .power_up = "low";

cycloneive_lcell_comb \mem~296 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~204_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~140_q ),
	.cin(gnd),
	.combout(\mem~296_combout ),
	.cout());
defparam \mem~296 .lut_mask = 16'hFFDE;
defparam \mem~296 .sum_lutc_input = "datac";

dffeas \mem~236 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~236_q ),
	.prn(vcc));
defparam \mem~236 .is_wysiwyg = "true";
defparam \mem~236 .power_up = "low";

cycloneive_lcell_comb \mem~297 (
	.dataa(\mem~172_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~296_combout ),
	.datad(\mem~236_q ),
	.cin(gnd),
	.combout(\mem~297_combout ),
	.cout());
defparam \mem~297 .lut_mask = 16'hFFBE;
defparam \mem~297 .sum_lutc_input = "datac";

dffeas \mem~76 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~76_q ),
	.prn(vcc));
defparam \mem~76 .is_wysiwyg = "true";
defparam \mem~76 .power_up = "low";

dffeas \mem~44 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~44_q ),
	.prn(vcc));
defparam \mem~44 .is_wysiwyg = "true";
defparam \mem~44 .power_up = "low";

dffeas \mem~12 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~12_q ),
	.prn(vcc));
defparam \mem~12 .is_wysiwyg = "true";
defparam \mem~12 .power_up = "low";

cycloneive_lcell_comb \mem~298 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~44_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~12_q ),
	.cin(gnd),
	.combout(\mem~298_combout ),
	.cout());
defparam \mem~298 .lut_mask = 16'hFFDE;
defparam \mem~298 .sum_lutc_input = "datac";

dffeas \mem~108 (
	.clk(clk),
	.d(za_data_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~108_q ),
	.prn(vcc));
defparam \mem~108 .is_wysiwyg = "true";
defparam \mem~108 .power_up = "low";

cycloneive_lcell_comb \mem~299 (
	.dataa(\mem~76_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~298_combout ),
	.datad(\mem~108_q ),
	.cin(gnd),
	.combout(\mem~299_combout ),
	.cout());
defparam \mem~299 .lut_mask = 16'hFFBE;
defparam \mem~299 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~300 (
	.dataa(\mem~297_combout ),
	.datab(\mem~299_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~300_combout ),
	.cout());
defparam \mem~300 .lut_mask = 16'hAACC;
defparam \mem~300 .sum_lutc_input = "datac";

dffeas \internal_out_payload[12] (
	.clk(clk),
	.d(\mem~300_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[12]~q ),
	.prn(vcc));
defparam \internal_out_payload[12] .is_wysiwyg = "true";
defparam \internal_out_payload[12] .power_up = "low";

dffeas \mem~165 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~165_q ),
	.prn(vcc));
defparam \mem~165 .is_wysiwyg = "true";
defparam \mem~165 .power_up = "low";

dffeas \mem~197 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~197_q ),
	.prn(vcc));
defparam \mem~197 .is_wysiwyg = "true";
defparam \mem~197 .power_up = "low";

dffeas \mem~133 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~133_q ),
	.prn(vcc));
defparam \mem~133 .is_wysiwyg = "true";
defparam \mem~133 .power_up = "low";

cycloneive_lcell_comb \mem~301 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~197_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~133_q ),
	.cin(gnd),
	.combout(\mem~301_combout ),
	.cout());
defparam \mem~301 .lut_mask = 16'hFFDE;
defparam \mem~301 .sum_lutc_input = "datac";

dffeas \mem~229 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~229_q ),
	.prn(vcc));
defparam \mem~229 .is_wysiwyg = "true";
defparam \mem~229 .power_up = "low";

cycloneive_lcell_comb \mem~302 (
	.dataa(\mem~165_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~301_combout ),
	.datad(\mem~229_q ),
	.cin(gnd),
	.combout(\mem~302_combout ),
	.cout());
defparam \mem~302 .lut_mask = 16'hFFBE;
defparam \mem~302 .sum_lutc_input = "datac";

dffeas \mem~69 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~69_q ),
	.prn(vcc));
defparam \mem~69 .is_wysiwyg = "true";
defparam \mem~69 .power_up = "low";

dffeas \mem~37 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~37_q ),
	.prn(vcc));
defparam \mem~37 .is_wysiwyg = "true";
defparam \mem~37 .power_up = "low";

dffeas \mem~5 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~5_q ),
	.prn(vcc));
defparam \mem~5 .is_wysiwyg = "true";
defparam \mem~5 .power_up = "low";

cycloneive_lcell_comb \mem~303 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~37_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~5_q ),
	.cin(gnd),
	.combout(\mem~303_combout ),
	.cout());
defparam \mem~303 .lut_mask = 16'hFFDE;
defparam \mem~303 .sum_lutc_input = "datac";

dffeas \mem~101 (
	.clk(clk),
	.d(za_data_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~101_q ),
	.prn(vcc));
defparam \mem~101 .is_wysiwyg = "true";
defparam \mem~101 .power_up = "low";

cycloneive_lcell_comb \mem~304 (
	.dataa(\mem~69_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~303_combout ),
	.datad(\mem~101_q ),
	.cin(gnd),
	.combout(\mem~304_combout ),
	.cout());
defparam \mem~304 .lut_mask = 16'hFFBE;
defparam \mem~304 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~305 (
	.dataa(\mem~302_combout ),
	.datab(\mem~304_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~305_combout ),
	.cout());
defparam \mem~305 .lut_mask = 16'hAACC;
defparam \mem~305 .sum_lutc_input = "datac";

dffeas \internal_out_payload[5] (
	.clk(clk),
	.d(\mem~305_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[5]~q ),
	.prn(vcc));
defparam \internal_out_payload[5] .is_wysiwyg = "true";
defparam \internal_out_payload[5] .power_up = "low";

dffeas \mem~174 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~174_q ),
	.prn(vcc));
defparam \mem~174 .is_wysiwyg = "true";
defparam \mem~174 .power_up = "low";

dffeas \mem~206 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~206_q ),
	.prn(vcc));
defparam \mem~206 .is_wysiwyg = "true";
defparam \mem~206 .power_up = "low";

dffeas \mem~142 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~142_q ),
	.prn(vcc));
defparam \mem~142 .is_wysiwyg = "true";
defparam \mem~142 .power_up = "low";

cycloneive_lcell_comb \mem~306 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~206_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~142_q ),
	.cin(gnd),
	.combout(\mem~306_combout ),
	.cout());
defparam \mem~306 .lut_mask = 16'hFFDE;
defparam \mem~306 .sum_lutc_input = "datac";

dffeas \mem~238 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~238_q ),
	.prn(vcc));
defparam \mem~238 .is_wysiwyg = "true";
defparam \mem~238 .power_up = "low";

cycloneive_lcell_comb \mem~307 (
	.dataa(\mem~174_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~306_combout ),
	.datad(\mem~238_q ),
	.cin(gnd),
	.combout(\mem~307_combout ),
	.cout());
defparam \mem~307 .lut_mask = 16'hFFBE;
defparam \mem~307 .sum_lutc_input = "datac";

dffeas \mem~78 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~78_q ),
	.prn(vcc));
defparam \mem~78 .is_wysiwyg = "true";
defparam \mem~78 .power_up = "low";

dffeas \mem~46 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~46_q ),
	.prn(vcc));
defparam \mem~46 .is_wysiwyg = "true";
defparam \mem~46 .power_up = "low";

dffeas \mem~14 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~14_q ),
	.prn(vcc));
defparam \mem~14 .is_wysiwyg = "true";
defparam \mem~14 .power_up = "low";

cycloneive_lcell_comb \mem~308 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~46_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~14_q ),
	.cin(gnd),
	.combout(\mem~308_combout ),
	.cout());
defparam \mem~308 .lut_mask = 16'hFFDE;
defparam \mem~308 .sum_lutc_input = "datac";

dffeas \mem~110 (
	.clk(clk),
	.d(za_data_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~110_q ),
	.prn(vcc));
defparam \mem~110 .is_wysiwyg = "true";
defparam \mem~110 .power_up = "low";

cycloneive_lcell_comb \mem~309 (
	.dataa(\mem~78_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~308_combout ),
	.datad(\mem~110_q ),
	.cin(gnd),
	.combout(\mem~309_combout ),
	.cout());
defparam \mem~309 .lut_mask = 16'hFFBE;
defparam \mem~309 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~310 (
	.dataa(\mem~307_combout ),
	.datab(\mem~309_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~310_combout ),
	.cout());
defparam \mem~310 .lut_mask = 16'hAACC;
defparam \mem~310 .sum_lutc_input = "datac";

dffeas \internal_out_payload[14] (
	.clk(clk),
	.d(\mem~310_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[14]~q ),
	.prn(vcc));
defparam \internal_out_payload[14] .is_wysiwyg = "true";
defparam \internal_out_payload[14] .power_up = "low";

dffeas \mem~175 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~175_q ),
	.prn(vcc));
defparam \mem~175 .is_wysiwyg = "true";
defparam \mem~175 .power_up = "low";

dffeas \mem~207 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~207_q ),
	.prn(vcc));
defparam \mem~207 .is_wysiwyg = "true";
defparam \mem~207 .power_up = "low";

dffeas \mem~143 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~143_q ),
	.prn(vcc));
defparam \mem~143 .is_wysiwyg = "true";
defparam \mem~143 .power_up = "low";

cycloneive_lcell_comb \mem~311 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~207_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~143_q ),
	.cin(gnd),
	.combout(\mem~311_combout ),
	.cout());
defparam \mem~311 .lut_mask = 16'hFFDE;
defparam \mem~311 .sum_lutc_input = "datac";

dffeas \mem~239 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~239_q ),
	.prn(vcc));
defparam \mem~239 .is_wysiwyg = "true";
defparam \mem~239 .power_up = "low";

cycloneive_lcell_comb \mem~312 (
	.dataa(\mem~175_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~311_combout ),
	.datad(\mem~239_q ),
	.cin(gnd),
	.combout(\mem~312_combout ),
	.cout());
defparam \mem~312 .lut_mask = 16'hFFBE;
defparam \mem~312 .sum_lutc_input = "datac";

dffeas \mem~79 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~79_q ),
	.prn(vcc));
defparam \mem~79 .is_wysiwyg = "true";
defparam \mem~79 .power_up = "low";

dffeas \mem~47 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~47_q ),
	.prn(vcc));
defparam \mem~47 .is_wysiwyg = "true";
defparam \mem~47 .power_up = "low";

dffeas \mem~15 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~15_q ),
	.prn(vcc));
defparam \mem~15 .is_wysiwyg = "true";
defparam \mem~15 .power_up = "low";

cycloneive_lcell_comb \mem~313 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~47_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~15_q ),
	.cin(gnd),
	.combout(\mem~313_combout ),
	.cout());
defparam \mem~313 .lut_mask = 16'hFFDE;
defparam \mem~313 .sum_lutc_input = "datac";

dffeas \mem~111 (
	.clk(clk),
	.d(za_data_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~111_q ),
	.prn(vcc));
defparam \mem~111 .is_wysiwyg = "true";
defparam \mem~111 .power_up = "low";

cycloneive_lcell_comb \mem~314 (
	.dataa(\mem~79_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~313_combout ),
	.datad(\mem~111_q ),
	.cin(gnd),
	.combout(\mem~314_combout ),
	.cout());
defparam \mem~314 .lut_mask = 16'hFFBE;
defparam \mem~314 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~315 (
	.dataa(\mem~312_combout ),
	.datab(\mem~314_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~315_combout ),
	.cout());
defparam \mem~315 .lut_mask = 16'hAACC;
defparam \mem~315 .sum_lutc_input = "datac";

dffeas \internal_out_payload[15] (
	.clk(clk),
	.d(\mem~315_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[15]~q ),
	.prn(vcc));
defparam \internal_out_payload[15] .is_wysiwyg = "true";
defparam \internal_out_payload[15] .power_up = "low";

dffeas \mem~181 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~181_q ),
	.prn(vcc));
defparam \mem~181 .is_wysiwyg = "true";
defparam \mem~181 .power_up = "low";

dffeas \mem~213 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~213_q ),
	.prn(vcc));
defparam \mem~213 .is_wysiwyg = "true";
defparam \mem~213 .power_up = "low";

dffeas \mem~149 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~149_q ),
	.prn(vcc));
defparam \mem~149 .is_wysiwyg = "true";
defparam \mem~149 .power_up = "low";

cycloneive_lcell_comb \mem~316 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~213_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~149_q ),
	.cin(gnd),
	.combout(\mem~316_combout ),
	.cout());
defparam \mem~316 .lut_mask = 16'hFFDE;
defparam \mem~316 .sum_lutc_input = "datac";

dffeas \mem~245 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~245_q ),
	.prn(vcc));
defparam \mem~245 .is_wysiwyg = "true";
defparam \mem~245 .power_up = "low";

cycloneive_lcell_comb \mem~317 (
	.dataa(\mem~181_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~316_combout ),
	.datad(\mem~245_q ),
	.cin(gnd),
	.combout(\mem~317_combout ),
	.cout());
defparam \mem~317 .lut_mask = 16'hFFBE;
defparam \mem~317 .sum_lutc_input = "datac";

dffeas \mem~85 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~85_q ),
	.prn(vcc));
defparam \mem~85 .is_wysiwyg = "true";
defparam \mem~85 .power_up = "low";

dffeas \mem~53 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~53_q ),
	.prn(vcc));
defparam \mem~53 .is_wysiwyg = "true";
defparam \mem~53 .power_up = "low";

dffeas \mem~21 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~21_q ),
	.prn(vcc));
defparam \mem~21 .is_wysiwyg = "true";
defparam \mem~21 .power_up = "low";

cycloneive_lcell_comb \mem~318 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~53_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~21_q ),
	.cin(gnd),
	.combout(\mem~318_combout ),
	.cout());
defparam \mem~318 .lut_mask = 16'hFFDE;
defparam \mem~318 .sum_lutc_input = "datac";

dffeas \mem~117 (
	.clk(clk),
	.d(za_data_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~117_q ),
	.prn(vcc));
defparam \mem~117 .is_wysiwyg = "true";
defparam \mem~117 .power_up = "low";

cycloneive_lcell_comb \mem~319 (
	.dataa(\mem~85_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~318_combout ),
	.datad(\mem~117_q ),
	.cin(gnd),
	.combout(\mem~319_combout ),
	.cout());
defparam \mem~319 .lut_mask = 16'hFFBE;
defparam \mem~319 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~320 (
	.dataa(\mem~317_combout ),
	.datab(\mem~319_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~320_combout ),
	.cout());
defparam \mem~320 .lut_mask = 16'hAACC;
defparam \mem~320 .sum_lutc_input = "datac";

dffeas \internal_out_payload[21] (
	.clk(clk),
	.d(\mem~320_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[21]~q ),
	.prn(vcc));
defparam \internal_out_payload[21] .is_wysiwyg = "true";
defparam \internal_out_payload[21] .power_up = "low";

dffeas \mem~178 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~178_q ),
	.prn(vcc));
defparam \mem~178 .is_wysiwyg = "true";
defparam \mem~178 .power_up = "low";

dffeas \mem~210 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~210_q ),
	.prn(vcc));
defparam \mem~210 .is_wysiwyg = "true";
defparam \mem~210 .power_up = "low";

dffeas \mem~146 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~146_q ),
	.prn(vcc));
defparam \mem~146 .is_wysiwyg = "true";
defparam \mem~146 .power_up = "low";

cycloneive_lcell_comb \mem~321 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~210_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~146_q ),
	.cin(gnd),
	.combout(\mem~321_combout ),
	.cout());
defparam \mem~321 .lut_mask = 16'hFFDE;
defparam \mem~321 .sum_lutc_input = "datac";

dffeas \mem~242 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~242_q ),
	.prn(vcc));
defparam \mem~242 .is_wysiwyg = "true";
defparam \mem~242 .power_up = "low";

cycloneive_lcell_comb \mem~322 (
	.dataa(\mem~178_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~321_combout ),
	.datad(\mem~242_q ),
	.cin(gnd),
	.combout(\mem~322_combout ),
	.cout());
defparam \mem~322 .lut_mask = 16'hFFBE;
defparam \mem~322 .sum_lutc_input = "datac";

dffeas \mem~82 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~82_q ),
	.prn(vcc));
defparam \mem~82 .is_wysiwyg = "true";
defparam \mem~82 .power_up = "low";

dffeas \mem~50 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~50_q ),
	.prn(vcc));
defparam \mem~50 .is_wysiwyg = "true";
defparam \mem~50 .power_up = "low";

dffeas \mem~18 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~18_q ),
	.prn(vcc));
defparam \mem~18 .is_wysiwyg = "true";
defparam \mem~18 .power_up = "low";

cycloneive_lcell_comb \mem~323 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~50_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~18_q ),
	.cin(gnd),
	.combout(\mem~323_combout ),
	.cout());
defparam \mem~323 .lut_mask = 16'hFFDE;
defparam \mem~323 .sum_lutc_input = "datac";

dffeas \mem~114 (
	.clk(clk),
	.d(za_data_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~114_q ),
	.prn(vcc));
defparam \mem~114 .is_wysiwyg = "true";
defparam \mem~114 .power_up = "low";

cycloneive_lcell_comb \mem~324 (
	.dataa(\mem~82_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~323_combout ),
	.datad(\mem~114_q ),
	.cin(gnd),
	.combout(\mem~324_combout ),
	.cout());
defparam \mem~324 .lut_mask = 16'hFFBE;
defparam \mem~324 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~325 (
	.dataa(\mem~322_combout ),
	.datab(\mem~324_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~325_combout ),
	.cout());
defparam \mem~325 .lut_mask = 16'hAACC;
defparam \mem~325 .sum_lutc_input = "datac";

dffeas \internal_out_payload[18] (
	.clk(clk),
	.d(\mem~325_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[18]~q ),
	.prn(vcc));
defparam \internal_out_payload[18] .is_wysiwyg = "true";
defparam \internal_out_payload[18] .power_up = "low";

dffeas \mem~177 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~177_q ),
	.prn(vcc));
defparam \mem~177 .is_wysiwyg = "true";
defparam \mem~177 .power_up = "low";

dffeas \mem~209 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~209_q ),
	.prn(vcc));
defparam \mem~209 .is_wysiwyg = "true";
defparam \mem~209 .power_up = "low";

dffeas \mem~145 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~145_q ),
	.prn(vcc));
defparam \mem~145 .is_wysiwyg = "true";
defparam \mem~145 .power_up = "low";

cycloneive_lcell_comb \mem~326 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~209_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~145_q ),
	.cin(gnd),
	.combout(\mem~326_combout ),
	.cout());
defparam \mem~326 .lut_mask = 16'hFFDE;
defparam \mem~326 .sum_lutc_input = "datac";

dffeas \mem~241 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~241_q ),
	.prn(vcc));
defparam \mem~241 .is_wysiwyg = "true";
defparam \mem~241 .power_up = "low";

cycloneive_lcell_comb \mem~327 (
	.dataa(\mem~177_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~326_combout ),
	.datad(\mem~241_q ),
	.cin(gnd),
	.combout(\mem~327_combout ),
	.cout());
defparam \mem~327 .lut_mask = 16'hFFBE;
defparam \mem~327 .sum_lutc_input = "datac";

dffeas \mem~81 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~81_q ),
	.prn(vcc));
defparam \mem~81 .is_wysiwyg = "true";
defparam \mem~81 .power_up = "low";

dffeas \mem~49 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~49_q ),
	.prn(vcc));
defparam \mem~49 .is_wysiwyg = "true";
defparam \mem~49 .power_up = "low";

dffeas \mem~17 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~17_q ),
	.prn(vcc));
defparam \mem~17 .is_wysiwyg = "true";
defparam \mem~17 .power_up = "low";

cycloneive_lcell_comb \mem~328 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~49_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~17_q ),
	.cin(gnd),
	.combout(\mem~328_combout ),
	.cout());
defparam \mem~328 .lut_mask = 16'hFFDE;
defparam \mem~328 .sum_lutc_input = "datac";

dffeas \mem~113 (
	.clk(clk),
	.d(za_data_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~113_q ),
	.prn(vcc));
defparam \mem~113 .is_wysiwyg = "true";
defparam \mem~113 .power_up = "low";

cycloneive_lcell_comb \mem~329 (
	.dataa(\mem~81_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~328_combout ),
	.datad(\mem~113_q ),
	.cin(gnd),
	.combout(\mem~329_combout ),
	.cout());
defparam \mem~329 .lut_mask = 16'hFFBE;
defparam \mem~329 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~330 (
	.dataa(\mem~327_combout ),
	.datab(\mem~329_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~330_combout ),
	.cout());
defparam \mem~330 .lut_mask = 16'hAACC;
defparam \mem~330 .sum_lutc_input = "datac";

dffeas \internal_out_payload[17] (
	.clk(clk),
	.d(\mem~330_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[17]~q ),
	.prn(vcc));
defparam \internal_out_payload[17] .is_wysiwyg = "true";
defparam \internal_out_payload[17] .power_up = "low";

dffeas \mem~191 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~191_q ),
	.prn(vcc));
defparam \mem~191 .is_wysiwyg = "true";
defparam \mem~191 .power_up = "low";

dffeas \mem~223 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~223_q ),
	.prn(vcc));
defparam \mem~223 .is_wysiwyg = "true";
defparam \mem~223 .power_up = "low";

dffeas \mem~159 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~159_q ),
	.prn(vcc));
defparam \mem~159 .is_wysiwyg = "true";
defparam \mem~159 .power_up = "low";

cycloneive_lcell_comb \mem~331 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~223_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~159_q ),
	.cin(gnd),
	.combout(\mem~331_combout ),
	.cout());
defparam \mem~331 .lut_mask = 16'hFFDE;
defparam \mem~331 .sum_lutc_input = "datac";

dffeas \mem~255 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~255_q ),
	.prn(vcc));
defparam \mem~255 .is_wysiwyg = "true";
defparam \mem~255 .power_up = "low";

cycloneive_lcell_comb \mem~332 (
	.dataa(\mem~191_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~331_combout ),
	.datad(\mem~255_q ),
	.cin(gnd),
	.combout(\mem~332_combout ),
	.cout());
defparam \mem~332 .lut_mask = 16'hFFBE;
defparam \mem~332 .sum_lutc_input = "datac";

dffeas \mem~95 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~95_q ),
	.prn(vcc));
defparam \mem~95 .is_wysiwyg = "true";
defparam \mem~95 .power_up = "low";

dffeas \mem~63 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~63_q ),
	.prn(vcc));
defparam \mem~63 .is_wysiwyg = "true";
defparam \mem~63 .power_up = "low";

dffeas \mem~31 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~31_q ),
	.prn(vcc));
defparam \mem~31 .is_wysiwyg = "true";
defparam \mem~31 .power_up = "low";

cycloneive_lcell_comb \mem~333 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~63_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~31_q ),
	.cin(gnd),
	.combout(\mem~333_combout ),
	.cout());
defparam \mem~333 .lut_mask = 16'hFFDE;
defparam \mem~333 .sum_lutc_input = "datac";

dffeas \mem~127 (
	.clk(clk),
	.d(za_data_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~127_q ),
	.prn(vcc));
defparam \mem~127 .is_wysiwyg = "true";
defparam \mem~127 .power_up = "low";

cycloneive_lcell_comb \mem~334 (
	.dataa(\mem~95_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~333_combout ),
	.datad(\mem~127_q ),
	.cin(gnd),
	.combout(\mem~334_combout ),
	.cout());
defparam \mem~334 .lut_mask = 16'hFFBE;
defparam \mem~334 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~335 (
	.dataa(\mem~332_combout ),
	.datab(\mem~334_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~335_combout ),
	.cout());
defparam \mem~335 .lut_mask = 16'hAACC;
defparam \mem~335 .sum_lutc_input = "datac";

dffeas \internal_out_payload[31] (
	.clk(clk),
	.d(\mem~335_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[31]~q ),
	.prn(vcc));
defparam \internal_out_payload[31] .is_wysiwyg = "true";
defparam \internal_out_payload[31] .power_up = "low";

dffeas \mem~190 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~190_q ),
	.prn(vcc));
defparam \mem~190 .is_wysiwyg = "true";
defparam \mem~190 .power_up = "low";

dffeas \mem~222 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~222_q ),
	.prn(vcc));
defparam \mem~222 .is_wysiwyg = "true";
defparam \mem~222 .power_up = "low";

dffeas \mem~158 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~158_q ),
	.prn(vcc));
defparam \mem~158 .is_wysiwyg = "true";
defparam \mem~158 .power_up = "low";

cycloneive_lcell_comb \mem~336 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~222_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~158_q ),
	.cin(gnd),
	.combout(\mem~336_combout ),
	.cout());
defparam \mem~336 .lut_mask = 16'hFFDE;
defparam \mem~336 .sum_lutc_input = "datac";

dffeas \mem~254 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~254_q ),
	.prn(vcc));
defparam \mem~254 .is_wysiwyg = "true";
defparam \mem~254 .power_up = "low";

cycloneive_lcell_comb \mem~337 (
	.dataa(\mem~190_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~336_combout ),
	.datad(\mem~254_q ),
	.cin(gnd),
	.combout(\mem~337_combout ),
	.cout());
defparam \mem~337 .lut_mask = 16'hFFBE;
defparam \mem~337 .sum_lutc_input = "datac";

dffeas \mem~94 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~94_q ),
	.prn(vcc));
defparam \mem~94 .is_wysiwyg = "true";
defparam \mem~94 .power_up = "low";

dffeas \mem~62 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~62_q ),
	.prn(vcc));
defparam \mem~62 .is_wysiwyg = "true";
defparam \mem~62 .power_up = "low";

dffeas \mem~30 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~30_q ),
	.prn(vcc));
defparam \mem~30 .is_wysiwyg = "true";
defparam \mem~30 .power_up = "low";

cycloneive_lcell_comb \mem~338 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~62_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~30_q ),
	.cin(gnd),
	.combout(\mem~338_combout ),
	.cout());
defparam \mem~338 .lut_mask = 16'hFFDE;
defparam \mem~338 .sum_lutc_input = "datac";

dffeas \mem~126 (
	.clk(clk),
	.d(za_data_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~126_q ),
	.prn(vcc));
defparam \mem~126 .is_wysiwyg = "true";
defparam \mem~126 .power_up = "low";

cycloneive_lcell_comb \mem~339 (
	.dataa(\mem~94_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~338_combout ),
	.datad(\mem~126_q ),
	.cin(gnd),
	.combout(\mem~339_combout ),
	.cout());
defparam \mem~339 .lut_mask = 16'hFFBE;
defparam \mem~339 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~340 (
	.dataa(\mem~337_combout ),
	.datab(\mem~339_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~340_combout ),
	.cout());
defparam \mem~340 .lut_mask = 16'hAACC;
defparam \mem~340 .sum_lutc_input = "datac";

dffeas \internal_out_payload[30] (
	.clk(clk),
	.d(\mem~340_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[30]~q ),
	.prn(vcc));
defparam \internal_out_payload[30] .is_wysiwyg = "true";
defparam \internal_out_payload[30] .power_up = "low";

dffeas \mem~189 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~189_q ),
	.prn(vcc));
defparam \mem~189 .is_wysiwyg = "true";
defparam \mem~189 .power_up = "low";

dffeas \mem~221 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~221_q ),
	.prn(vcc));
defparam \mem~221 .is_wysiwyg = "true";
defparam \mem~221 .power_up = "low";

dffeas \mem~157 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~157_q ),
	.prn(vcc));
defparam \mem~157 .is_wysiwyg = "true";
defparam \mem~157 .power_up = "low";

cycloneive_lcell_comb \mem~341 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~221_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~157_q ),
	.cin(gnd),
	.combout(\mem~341_combout ),
	.cout());
defparam \mem~341 .lut_mask = 16'hFFDE;
defparam \mem~341 .sum_lutc_input = "datac";

dffeas \mem~253 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~253_q ),
	.prn(vcc));
defparam \mem~253 .is_wysiwyg = "true";
defparam \mem~253 .power_up = "low";

cycloneive_lcell_comb \mem~342 (
	.dataa(\mem~189_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~341_combout ),
	.datad(\mem~253_q ),
	.cin(gnd),
	.combout(\mem~342_combout ),
	.cout());
defparam \mem~342 .lut_mask = 16'hFFBE;
defparam \mem~342 .sum_lutc_input = "datac";

dffeas \mem~93 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~93_q ),
	.prn(vcc));
defparam \mem~93 .is_wysiwyg = "true";
defparam \mem~93 .power_up = "low";

dffeas \mem~61 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~61_q ),
	.prn(vcc));
defparam \mem~61 .is_wysiwyg = "true";
defparam \mem~61 .power_up = "low";

dffeas \mem~29 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~29_q ),
	.prn(vcc));
defparam \mem~29 .is_wysiwyg = "true";
defparam \mem~29 .power_up = "low";

cycloneive_lcell_comb \mem~343 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~61_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~29_q ),
	.cin(gnd),
	.combout(\mem~343_combout ),
	.cout());
defparam \mem~343 .lut_mask = 16'hFFDE;
defparam \mem~343 .sum_lutc_input = "datac";

dffeas \mem~125 (
	.clk(clk),
	.d(za_data_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~125_q ),
	.prn(vcc));
defparam \mem~125 .is_wysiwyg = "true";
defparam \mem~125 .power_up = "low";

cycloneive_lcell_comb \mem~344 (
	.dataa(\mem~93_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~343_combout ),
	.datad(\mem~125_q ),
	.cin(gnd),
	.combout(\mem~344_combout ),
	.cout());
defparam \mem~344 .lut_mask = 16'hFFBE;
defparam \mem~344 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~345 (
	.dataa(\mem~342_combout ),
	.datab(\mem~344_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~345_combout ),
	.cout());
defparam \mem~345 .lut_mask = 16'hAACC;
defparam \mem~345 .sum_lutc_input = "datac";

dffeas \internal_out_payload[29] (
	.clk(clk),
	.d(\mem~345_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[29]~q ),
	.prn(vcc));
defparam \internal_out_payload[29] .is_wysiwyg = "true";
defparam \internal_out_payload[29] .power_up = "low";

dffeas \mem~188 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~188_q ),
	.prn(vcc));
defparam \mem~188 .is_wysiwyg = "true";
defparam \mem~188 .power_up = "low";

dffeas \mem~220 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~220_q ),
	.prn(vcc));
defparam \mem~220 .is_wysiwyg = "true";
defparam \mem~220 .power_up = "low";

dffeas \mem~156 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~156_q ),
	.prn(vcc));
defparam \mem~156 .is_wysiwyg = "true";
defparam \mem~156 .power_up = "low";

cycloneive_lcell_comb \mem~346 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~220_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~156_q ),
	.cin(gnd),
	.combout(\mem~346_combout ),
	.cout());
defparam \mem~346 .lut_mask = 16'hFFDE;
defparam \mem~346 .sum_lutc_input = "datac";

dffeas \mem~252 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~252_q ),
	.prn(vcc));
defparam \mem~252 .is_wysiwyg = "true";
defparam \mem~252 .power_up = "low";

cycloneive_lcell_comb \mem~347 (
	.dataa(\mem~188_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~346_combout ),
	.datad(\mem~252_q ),
	.cin(gnd),
	.combout(\mem~347_combout ),
	.cout());
defparam \mem~347 .lut_mask = 16'hFFBE;
defparam \mem~347 .sum_lutc_input = "datac";

dffeas \mem~92 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~92_q ),
	.prn(vcc));
defparam \mem~92 .is_wysiwyg = "true";
defparam \mem~92 .power_up = "low";

dffeas \mem~60 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~60_q ),
	.prn(vcc));
defparam \mem~60 .is_wysiwyg = "true";
defparam \mem~60 .power_up = "low";

dffeas \mem~28 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~28_q ),
	.prn(vcc));
defparam \mem~28 .is_wysiwyg = "true";
defparam \mem~28 .power_up = "low";

cycloneive_lcell_comb \mem~348 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~60_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~28_q ),
	.cin(gnd),
	.combout(\mem~348_combout ),
	.cout());
defparam \mem~348 .lut_mask = 16'hFFDE;
defparam \mem~348 .sum_lutc_input = "datac";

dffeas \mem~124 (
	.clk(clk),
	.d(za_data_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~124_q ),
	.prn(vcc));
defparam \mem~124 .is_wysiwyg = "true";
defparam \mem~124 .power_up = "low";

cycloneive_lcell_comb \mem~349 (
	.dataa(\mem~92_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~348_combout ),
	.datad(\mem~124_q ),
	.cin(gnd),
	.combout(\mem~349_combout ),
	.cout());
defparam \mem~349 .lut_mask = 16'hFFBE;
defparam \mem~349 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~350 (
	.dataa(\mem~347_combout ),
	.datab(\mem~349_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~350_combout ),
	.cout());
defparam \mem~350 .lut_mask = 16'hAACC;
defparam \mem~350 .sum_lutc_input = "datac";

dffeas \internal_out_payload[28] (
	.clk(clk),
	.d(\mem~350_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[28]~q ),
	.prn(vcc));
defparam \internal_out_payload[28] .is_wysiwyg = "true";
defparam \internal_out_payload[28] .power_up = "low";

dffeas \mem~187 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~187_q ),
	.prn(vcc));
defparam \mem~187 .is_wysiwyg = "true";
defparam \mem~187 .power_up = "low";

dffeas \mem~219 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~219_q ),
	.prn(vcc));
defparam \mem~219 .is_wysiwyg = "true";
defparam \mem~219 .power_up = "low";

dffeas \mem~155 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~155_q ),
	.prn(vcc));
defparam \mem~155 .is_wysiwyg = "true";
defparam \mem~155 .power_up = "low";

cycloneive_lcell_comb \mem~351 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~219_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~155_q ),
	.cin(gnd),
	.combout(\mem~351_combout ),
	.cout());
defparam \mem~351 .lut_mask = 16'hFFDE;
defparam \mem~351 .sum_lutc_input = "datac";

dffeas \mem~251 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~251_q ),
	.prn(vcc));
defparam \mem~251 .is_wysiwyg = "true";
defparam \mem~251 .power_up = "low";

cycloneive_lcell_comb \mem~352 (
	.dataa(\mem~187_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~351_combout ),
	.datad(\mem~251_q ),
	.cin(gnd),
	.combout(\mem~352_combout ),
	.cout());
defparam \mem~352 .lut_mask = 16'hFFBE;
defparam \mem~352 .sum_lutc_input = "datac";

dffeas \mem~91 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~91_q ),
	.prn(vcc));
defparam \mem~91 .is_wysiwyg = "true";
defparam \mem~91 .power_up = "low";

dffeas \mem~59 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~59_q ),
	.prn(vcc));
defparam \mem~59 .is_wysiwyg = "true";
defparam \mem~59 .power_up = "low";

dffeas \mem~27 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~27_q ),
	.prn(vcc));
defparam \mem~27 .is_wysiwyg = "true";
defparam \mem~27 .power_up = "low";

cycloneive_lcell_comb \mem~353 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~59_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~27_q ),
	.cin(gnd),
	.combout(\mem~353_combout ),
	.cout());
defparam \mem~353 .lut_mask = 16'hFFDE;
defparam \mem~353 .sum_lutc_input = "datac";

dffeas \mem~123 (
	.clk(clk),
	.d(za_data_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~123_q ),
	.prn(vcc));
defparam \mem~123 .is_wysiwyg = "true";
defparam \mem~123 .power_up = "low";

cycloneive_lcell_comb \mem~354 (
	.dataa(\mem~91_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~353_combout ),
	.datad(\mem~123_q ),
	.cin(gnd),
	.combout(\mem~354_combout ),
	.cout());
defparam \mem~354 .lut_mask = 16'hFFBE;
defparam \mem~354 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~355 (
	.dataa(\mem~352_combout ),
	.datab(\mem~354_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~355_combout ),
	.cout());
defparam \mem~355 .lut_mask = 16'hAACC;
defparam \mem~355 .sum_lutc_input = "datac";

dffeas \internal_out_payload[27] (
	.clk(clk),
	.d(\mem~355_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[27]~q ),
	.prn(vcc));
defparam \internal_out_payload[27] .is_wysiwyg = "true";
defparam \internal_out_payload[27] .power_up = "low";

dffeas \mem~186 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~186_q ),
	.prn(vcc));
defparam \mem~186 .is_wysiwyg = "true";
defparam \mem~186 .power_up = "low";

dffeas \mem~218 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~218_q ),
	.prn(vcc));
defparam \mem~218 .is_wysiwyg = "true";
defparam \mem~218 .power_up = "low";

dffeas \mem~154 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~154_q ),
	.prn(vcc));
defparam \mem~154 .is_wysiwyg = "true";
defparam \mem~154 .power_up = "low";

cycloneive_lcell_comb \mem~356 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~218_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~154_q ),
	.cin(gnd),
	.combout(\mem~356_combout ),
	.cout());
defparam \mem~356 .lut_mask = 16'hFFDE;
defparam \mem~356 .sum_lutc_input = "datac";

dffeas \mem~250 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~250_q ),
	.prn(vcc));
defparam \mem~250 .is_wysiwyg = "true";
defparam \mem~250 .power_up = "low";

cycloneive_lcell_comb \mem~357 (
	.dataa(\mem~186_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~356_combout ),
	.datad(\mem~250_q ),
	.cin(gnd),
	.combout(\mem~357_combout ),
	.cout());
defparam \mem~357 .lut_mask = 16'hFFBE;
defparam \mem~357 .sum_lutc_input = "datac";

dffeas \mem~90 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~90_q ),
	.prn(vcc));
defparam \mem~90 .is_wysiwyg = "true";
defparam \mem~90 .power_up = "low";

dffeas \mem~58 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~58_q ),
	.prn(vcc));
defparam \mem~58 .is_wysiwyg = "true";
defparam \mem~58 .power_up = "low";

dffeas \mem~26 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~26_q ),
	.prn(vcc));
defparam \mem~26 .is_wysiwyg = "true";
defparam \mem~26 .power_up = "low";

cycloneive_lcell_comb \mem~358 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~58_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~26_q ),
	.cin(gnd),
	.combout(\mem~358_combout ),
	.cout());
defparam \mem~358 .lut_mask = 16'hFFDE;
defparam \mem~358 .sum_lutc_input = "datac";

dffeas \mem~122 (
	.clk(clk),
	.d(za_data_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~122_q ),
	.prn(vcc));
defparam \mem~122 .is_wysiwyg = "true";
defparam \mem~122 .power_up = "low";

cycloneive_lcell_comb \mem~359 (
	.dataa(\mem~90_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~358_combout ),
	.datad(\mem~122_q ),
	.cin(gnd),
	.combout(\mem~359_combout ),
	.cout());
defparam \mem~359 .lut_mask = 16'hFFBE;
defparam \mem~359 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~360 (
	.dataa(\mem~357_combout ),
	.datab(\mem~359_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~360_combout ),
	.cout());
defparam \mem~360 .lut_mask = 16'hAACC;
defparam \mem~360 .sum_lutc_input = "datac";

dffeas \internal_out_payload[26] (
	.clk(clk),
	.d(\mem~360_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[26]~q ),
	.prn(vcc));
defparam \internal_out_payload[26] .is_wysiwyg = "true";
defparam \internal_out_payload[26] .power_up = "low";

dffeas \mem~185 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~185_q ),
	.prn(vcc));
defparam \mem~185 .is_wysiwyg = "true";
defparam \mem~185 .power_up = "low";

dffeas \mem~217 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~217_q ),
	.prn(vcc));
defparam \mem~217 .is_wysiwyg = "true";
defparam \mem~217 .power_up = "low";

dffeas \mem~153 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~153_q ),
	.prn(vcc));
defparam \mem~153 .is_wysiwyg = "true";
defparam \mem~153 .power_up = "low";

cycloneive_lcell_comb \mem~361 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~217_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~153_q ),
	.cin(gnd),
	.combout(\mem~361_combout ),
	.cout());
defparam \mem~361 .lut_mask = 16'hFFDE;
defparam \mem~361 .sum_lutc_input = "datac";

dffeas \mem~249 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~249_q ),
	.prn(vcc));
defparam \mem~249 .is_wysiwyg = "true";
defparam \mem~249 .power_up = "low";

cycloneive_lcell_comb \mem~362 (
	.dataa(\mem~185_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~361_combout ),
	.datad(\mem~249_q ),
	.cin(gnd),
	.combout(\mem~362_combout ),
	.cout());
defparam \mem~362 .lut_mask = 16'hFFBE;
defparam \mem~362 .sum_lutc_input = "datac";

dffeas \mem~89 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~89_q ),
	.prn(vcc));
defparam \mem~89 .is_wysiwyg = "true";
defparam \mem~89 .power_up = "low";

dffeas \mem~57 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~57_q ),
	.prn(vcc));
defparam \mem~57 .is_wysiwyg = "true";
defparam \mem~57 .power_up = "low";

dffeas \mem~25 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~25_q ),
	.prn(vcc));
defparam \mem~25 .is_wysiwyg = "true";
defparam \mem~25 .power_up = "low";

cycloneive_lcell_comb \mem~363 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~57_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~25_q ),
	.cin(gnd),
	.combout(\mem~363_combout ),
	.cout());
defparam \mem~363 .lut_mask = 16'hFFDE;
defparam \mem~363 .sum_lutc_input = "datac";

dffeas \mem~121 (
	.clk(clk),
	.d(za_data_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~121_q ),
	.prn(vcc));
defparam \mem~121 .is_wysiwyg = "true";
defparam \mem~121 .power_up = "low";

cycloneive_lcell_comb \mem~364 (
	.dataa(\mem~89_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~363_combout ),
	.datad(\mem~121_q ),
	.cin(gnd),
	.combout(\mem~364_combout ),
	.cout());
defparam \mem~364 .lut_mask = 16'hFFBE;
defparam \mem~364 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~365 (
	.dataa(\mem~362_combout ),
	.datab(\mem~364_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~365_combout ),
	.cout());
defparam \mem~365 .lut_mask = 16'hAACC;
defparam \mem~365 .sum_lutc_input = "datac";

dffeas \internal_out_payload[25] (
	.clk(clk),
	.d(\mem~365_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[25]~q ),
	.prn(vcc));
defparam \internal_out_payload[25] .is_wysiwyg = "true";
defparam \internal_out_payload[25] .power_up = "low";

dffeas \mem~170 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~170_q ),
	.prn(vcc));
defparam \mem~170 .is_wysiwyg = "true";
defparam \mem~170 .power_up = "low";

dffeas \mem~202 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~202_q ),
	.prn(vcc));
defparam \mem~202 .is_wysiwyg = "true";
defparam \mem~202 .power_up = "low";

dffeas \mem~138 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~138_q ),
	.prn(vcc));
defparam \mem~138 .is_wysiwyg = "true";
defparam \mem~138 .power_up = "low";

cycloneive_lcell_comb \mem~366 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~202_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~138_q ),
	.cin(gnd),
	.combout(\mem~366_combout ),
	.cout());
defparam \mem~366 .lut_mask = 16'hFFDE;
defparam \mem~366 .sum_lutc_input = "datac";

dffeas \mem~234 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~234_q ),
	.prn(vcc));
defparam \mem~234 .is_wysiwyg = "true";
defparam \mem~234 .power_up = "low";

cycloneive_lcell_comb \mem~367 (
	.dataa(\mem~170_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~366_combout ),
	.datad(\mem~234_q ),
	.cin(gnd),
	.combout(\mem~367_combout ),
	.cout());
defparam \mem~367 .lut_mask = 16'hFFBE;
defparam \mem~367 .sum_lutc_input = "datac";

dffeas \mem~74 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~74_q ),
	.prn(vcc));
defparam \mem~74 .is_wysiwyg = "true";
defparam \mem~74 .power_up = "low";

dffeas \mem~42 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~42_q ),
	.prn(vcc));
defparam \mem~42 .is_wysiwyg = "true";
defparam \mem~42 .power_up = "low";

dffeas \mem~10 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~10_q ),
	.prn(vcc));
defparam \mem~10 .is_wysiwyg = "true";
defparam \mem~10 .power_up = "low";

cycloneive_lcell_comb \mem~368 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~42_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~10_q ),
	.cin(gnd),
	.combout(\mem~368_combout ),
	.cout());
defparam \mem~368 .lut_mask = 16'hFFDE;
defparam \mem~368 .sum_lutc_input = "datac";

dffeas \mem~106 (
	.clk(clk),
	.d(za_data_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~106_q ),
	.prn(vcc));
defparam \mem~106 .is_wysiwyg = "true";
defparam \mem~106 .power_up = "low";

cycloneive_lcell_comb \mem~369 (
	.dataa(\mem~74_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~368_combout ),
	.datad(\mem~106_q ),
	.cin(gnd),
	.combout(\mem~369_combout ),
	.cout());
defparam \mem~369 .lut_mask = 16'hFFBE;
defparam \mem~369 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~370 (
	.dataa(\mem~367_combout ),
	.datab(\mem~369_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~370_combout ),
	.cout());
defparam \mem~370 .lut_mask = 16'hAACC;
defparam \mem~370 .sum_lutc_input = "datac";

dffeas \internal_out_payload[10] (
	.clk(clk),
	.d(\mem~370_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[10]~q ),
	.prn(vcc));
defparam \internal_out_payload[10] .is_wysiwyg = "true";
defparam \internal_out_payload[10] .power_up = "low";

dffeas \mem~184 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~184_q ),
	.prn(vcc));
defparam \mem~184 .is_wysiwyg = "true";
defparam \mem~184 .power_up = "low";

dffeas \mem~216 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~216_q ),
	.prn(vcc));
defparam \mem~216 .is_wysiwyg = "true";
defparam \mem~216 .power_up = "low";

dffeas \mem~152 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~152_q ),
	.prn(vcc));
defparam \mem~152 .is_wysiwyg = "true";
defparam \mem~152 .power_up = "low";

cycloneive_lcell_comb \mem~371 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~216_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~152_q ),
	.cin(gnd),
	.combout(\mem~371_combout ),
	.cout());
defparam \mem~371 .lut_mask = 16'hFFDE;
defparam \mem~371 .sum_lutc_input = "datac";

dffeas \mem~248 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~248_q ),
	.prn(vcc));
defparam \mem~248 .is_wysiwyg = "true";
defparam \mem~248 .power_up = "low";

cycloneive_lcell_comb \mem~372 (
	.dataa(\mem~184_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~371_combout ),
	.datad(\mem~248_q ),
	.cin(gnd),
	.combout(\mem~372_combout ),
	.cout());
defparam \mem~372 .lut_mask = 16'hFFBE;
defparam \mem~372 .sum_lutc_input = "datac";

dffeas \mem~88 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~88_q ),
	.prn(vcc));
defparam \mem~88 .is_wysiwyg = "true";
defparam \mem~88 .power_up = "low";

dffeas \mem~56 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~56_q ),
	.prn(vcc));
defparam \mem~56 .is_wysiwyg = "true";
defparam \mem~56 .power_up = "low";

dffeas \mem~24 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~24_q ),
	.prn(vcc));
defparam \mem~24 .is_wysiwyg = "true";
defparam \mem~24 .power_up = "low";

cycloneive_lcell_comb \mem~373 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~56_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~24_q ),
	.cin(gnd),
	.combout(\mem~373_combout ),
	.cout());
defparam \mem~373 .lut_mask = 16'hFFDE;
defparam \mem~373 .sum_lutc_input = "datac";

dffeas \mem~120 (
	.clk(clk),
	.d(za_data_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~120_q ),
	.prn(vcc));
defparam \mem~120 .is_wysiwyg = "true";
defparam \mem~120 .power_up = "low";

cycloneive_lcell_comb \mem~374 (
	.dataa(\mem~88_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~373_combout ),
	.datad(\mem~120_q ),
	.cin(gnd),
	.combout(\mem~374_combout ),
	.cout());
defparam \mem~374 .lut_mask = 16'hFFBE;
defparam \mem~374 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~375 (
	.dataa(\mem~372_combout ),
	.datab(\mem~374_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~375_combout ),
	.cout());
defparam \mem~375 .lut_mask = 16'hAACC;
defparam \mem~375 .sum_lutc_input = "datac";

dffeas \internal_out_payload[24] (
	.clk(clk),
	.d(\mem~375_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[24]~q ),
	.prn(vcc));
defparam \internal_out_payload[24] .is_wysiwyg = "true";
defparam \internal_out_payload[24] .power_up = "low";

dffeas \mem~169 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~169_q ),
	.prn(vcc));
defparam \mem~169 .is_wysiwyg = "true";
defparam \mem~169 .power_up = "low";

dffeas \mem~201 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~201_q ),
	.prn(vcc));
defparam \mem~201 .is_wysiwyg = "true";
defparam \mem~201 .power_up = "low";

dffeas \mem~137 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~137_q ),
	.prn(vcc));
defparam \mem~137 .is_wysiwyg = "true";
defparam \mem~137 .power_up = "low";

cycloneive_lcell_comb \mem~376 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~201_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~137_q ),
	.cin(gnd),
	.combout(\mem~376_combout ),
	.cout());
defparam \mem~376 .lut_mask = 16'hFFDE;
defparam \mem~376 .sum_lutc_input = "datac";

dffeas \mem~233 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~233_q ),
	.prn(vcc));
defparam \mem~233 .is_wysiwyg = "true";
defparam \mem~233 .power_up = "low";

cycloneive_lcell_comb \mem~377 (
	.dataa(\mem~169_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~376_combout ),
	.datad(\mem~233_q ),
	.cin(gnd),
	.combout(\mem~377_combout ),
	.cout());
defparam \mem~377 .lut_mask = 16'hFFBE;
defparam \mem~377 .sum_lutc_input = "datac";

dffeas \mem~73 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~73_q ),
	.prn(vcc));
defparam \mem~73 .is_wysiwyg = "true";
defparam \mem~73 .power_up = "low";

dffeas \mem~41 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~41_q ),
	.prn(vcc));
defparam \mem~41 .is_wysiwyg = "true";
defparam \mem~41 .power_up = "low";

dffeas \mem~9 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~9_q ),
	.prn(vcc));
defparam \mem~9 .is_wysiwyg = "true";
defparam \mem~9 .power_up = "low";

cycloneive_lcell_comb \mem~378 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~41_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~9_q ),
	.cin(gnd),
	.combout(\mem~378_combout ),
	.cout());
defparam \mem~378 .lut_mask = 16'hFFDE;
defparam \mem~378 .sum_lutc_input = "datac";

dffeas \mem~105 (
	.clk(clk),
	.d(za_data_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~105_q ),
	.prn(vcc));
defparam \mem~105 .is_wysiwyg = "true";
defparam \mem~105 .power_up = "low";

cycloneive_lcell_comb \mem~379 (
	.dataa(\mem~73_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~378_combout ),
	.datad(\mem~105_q ),
	.cin(gnd),
	.combout(\mem~379_combout ),
	.cout());
defparam \mem~379 .lut_mask = 16'hFFBE;
defparam \mem~379 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~380 (
	.dataa(\mem~377_combout ),
	.datab(\mem~379_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~380_combout ),
	.cout());
defparam \mem~380 .lut_mask = 16'hAACC;
defparam \mem~380 .sum_lutc_input = "datac";

dffeas \internal_out_payload[9] (
	.clk(clk),
	.d(\mem~380_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[9]~q ),
	.prn(vcc));
defparam \internal_out_payload[9] .is_wysiwyg = "true";
defparam \internal_out_payload[9] .power_up = "low";

dffeas \mem~183 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~183_q ),
	.prn(vcc));
defparam \mem~183 .is_wysiwyg = "true";
defparam \mem~183 .power_up = "low";

dffeas \mem~215 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~215_q ),
	.prn(vcc));
defparam \mem~215 .is_wysiwyg = "true";
defparam \mem~215 .power_up = "low";

dffeas \mem~151 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~151_q ),
	.prn(vcc));
defparam \mem~151 .is_wysiwyg = "true";
defparam \mem~151 .power_up = "low";

cycloneive_lcell_comb \mem~381 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~215_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~151_q ),
	.cin(gnd),
	.combout(\mem~381_combout ),
	.cout());
defparam \mem~381 .lut_mask = 16'hFFDE;
defparam \mem~381 .sum_lutc_input = "datac";

dffeas \mem~247 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~247_q ),
	.prn(vcc));
defparam \mem~247 .is_wysiwyg = "true";
defparam \mem~247 .power_up = "low";

cycloneive_lcell_comb \mem~382 (
	.dataa(\mem~183_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~381_combout ),
	.datad(\mem~247_q ),
	.cin(gnd),
	.combout(\mem~382_combout ),
	.cout());
defparam \mem~382 .lut_mask = 16'hFFBE;
defparam \mem~382 .sum_lutc_input = "datac";

dffeas \mem~87 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~87_q ),
	.prn(vcc));
defparam \mem~87 .is_wysiwyg = "true";
defparam \mem~87 .power_up = "low";

dffeas \mem~55 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~55_q ),
	.prn(vcc));
defparam \mem~55 .is_wysiwyg = "true";
defparam \mem~55 .power_up = "low";

dffeas \mem~23 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~23_q ),
	.prn(vcc));
defparam \mem~23 .is_wysiwyg = "true";
defparam \mem~23 .power_up = "low";

cycloneive_lcell_comb \mem~383 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~55_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~23_q ),
	.cin(gnd),
	.combout(\mem~383_combout ),
	.cout());
defparam \mem~383 .lut_mask = 16'hFFDE;
defparam \mem~383 .sum_lutc_input = "datac";

dffeas \mem~119 (
	.clk(clk),
	.d(za_data_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~119_q ),
	.prn(vcc));
defparam \mem~119 .is_wysiwyg = "true";
defparam \mem~119 .power_up = "low";

cycloneive_lcell_comb \mem~384 (
	.dataa(\mem~87_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~383_combout ),
	.datad(\mem~119_q ),
	.cin(gnd),
	.combout(\mem~384_combout ),
	.cout());
defparam \mem~384 .lut_mask = 16'hFFBE;
defparam \mem~384 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~385 (
	.dataa(\mem~382_combout ),
	.datab(\mem~384_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~385_combout ),
	.cout());
defparam \mem~385 .lut_mask = 16'hAACC;
defparam \mem~385 .sum_lutc_input = "datac";

dffeas \internal_out_payload[23] (
	.clk(clk),
	.d(\mem~385_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[23]~q ),
	.prn(vcc));
defparam \internal_out_payload[23] .is_wysiwyg = "true";
defparam \internal_out_payload[23] .power_up = "low";

dffeas \mem~168 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~168_q ),
	.prn(vcc));
defparam \mem~168 .is_wysiwyg = "true";
defparam \mem~168 .power_up = "low";

dffeas \mem~200 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~200_q ),
	.prn(vcc));
defparam \mem~200 .is_wysiwyg = "true";
defparam \mem~200 .power_up = "low";

dffeas \mem~136 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~136_q ),
	.prn(vcc));
defparam \mem~136 .is_wysiwyg = "true";
defparam \mem~136 .power_up = "low";

cycloneive_lcell_comb \mem~386 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~200_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~136_q ),
	.cin(gnd),
	.combout(\mem~386_combout ),
	.cout());
defparam \mem~386 .lut_mask = 16'hFFDE;
defparam \mem~386 .sum_lutc_input = "datac";

dffeas \mem~232 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~232_q ),
	.prn(vcc));
defparam \mem~232 .is_wysiwyg = "true";
defparam \mem~232 .power_up = "low";

cycloneive_lcell_comb \mem~387 (
	.dataa(\mem~168_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~386_combout ),
	.datad(\mem~232_q ),
	.cin(gnd),
	.combout(\mem~387_combout ),
	.cout());
defparam \mem~387 .lut_mask = 16'hFFBE;
defparam \mem~387 .sum_lutc_input = "datac";

dffeas \mem~72 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~72_q ),
	.prn(vcc));
defparam \mem~72 .is_wysiwyg = "true";
defparam \mem~72 .power_up = "low";

dffeas \mem~40 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~40_q ),
	.prn(vcc));
defparam \mem~40 .is_wysiwyg = "true";
defparam \mem~40 .power_up = "low";

dffeas \mem~8 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~8_q ),
	.prn(vcc));
defparam \mem~8 .is_wysiwyg = "true";
defparam \mem~8 .power_up = "low";

cycloneive_lcell_comb \mem~388 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~40_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~8_q ),
	.cin(gnd),
	.combout(\mem~388_combout ),
	.cout());
defparam \mem~388 .lut_mask = 16'hFFDE;
defparam \mem~388 .sum_lutc_input = "datac";

dffeas \mem~104 (
	.clk(clk),
	.d(za_data_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~104_q ),
	.prn(vcc));
defparam \mem~104 .is_wysiwyg = "true";
defparam \mem~104 .power_up = "low";

cycloneive_lcell_comb \mem~389 (
	.dataa(\mem~72_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~388_combout ),
	.datad(\mem~104_q ),
	.cin(gnd),
	.combout(\mem~389_combout ),
	.cout());
defparam \mem~389 .lut_mask = 16'hFFBE;
defparam \mem~389 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~390 (
	.dataa(\mem~387_combout ),
	.datab(\mem~389_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~390_combout ),
	.cout());
defparam \mem~390 .lut_mask = 16'hAACC;
defparam \mem~390 .sum_lutc_input = "datac";

dffeas \internal_out_payload[8] (
	.clk(clk),
	.d(\mem~390_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[8]~q ),
	.prn(vcc));
defparam \internal_out_payload[8] .is_wysiwyg = "true";
defparam \internal_out_payload[8] .power_up = "low";

dffeas \mem~182 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~182_q ),
	.prn(vcc));
defparam \mem~182 .is_wysiwyg = "true";
defparam \mem~182 .power_up = "low";

dffeas \mem~214 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~214_q ),
	.prn(vcc));
defparam \mem~214 .is_wysiwyg = "true";
defparam \mem~214 .power_up = "low";

dffeas \mem~150 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~150_q ),
	.prn(vcc));
defparam \mem~150 .is_wysiwyg = "true";
defparam \mem~150 .power_up = "low";

cycloneive_lcell_comb \mem~391 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~214_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~150_q ),
	.cin(gnd),
	.combout(\mem~391_combout ),
	.cout());
defparam \mem~391 .lut_mask = 16'hFFDE;
defparam \mem~391 .sum_lutc_input = "datac";

dffeas \mem~246 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~246_q ),
	.prn(vcc));
defparam \mem~246 .is_wysiwyg = "true";
defparam \mem~246 .power_up = "low";

cycloneive_lcell_comb \mem~392 (
	.dataa(\mem~182_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~391_combout ),
	.datad(\mem~246_q ),
	.cin(gnd),
	.combout(\mem~392_combout ),
	.cout());
defparam \mem~392 .lut_mask = 16'hFFBE;
defparam \mem~392 .sum_lutc_input = "datac";

dffeas \mem~86 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~86_q ),
	.prn(vcc));
defparam \mem~86 .is_wysiwyg = "true";
defparam \mem~86 .power_up = "low";

dffeas \mem~54 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~54_q ),
	.prn(vcc));
defparam \mem~54 .is_wysiwyg = "true";
defparam \mem~54 .power_up = "low";

dffeas \mem~22 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~22_q ),
	.prn(vcc));
defparam \mem~22 .is_wysiwyg = "true";
defparam \mem~22 .power_up = "low";

cycloneive_lcell_comb \mem~393 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~54_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~22_q ),
	.cin(gnd),
	.combout(\mem~393_combout ),
	.cout());
defparam \mem~393 .lut_mask = 16'hFFDE;
defparam \mem~393 .sum_lutc_input = "datac";

dffeas \mem~118 (
	.clk(clk),
	.d(za_data_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~118_q ),
	.prn(vcc));
defparam \mem~118 .is_wysiwyg = "true";
defparam \mem~118 .power_up = "low";

cycloneive_lcell_comb \mem~394 (
	.dataa(\mem~86_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~393_combout ),
	.datad(\mem~118_q ),
	.cin(gnd),
	.combout(\mem~394_combout ),
	.cout());
defparam \mem~394 .lut_mask = 16'hFFBE;
defparam \mem~394 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~395 (
	.dataa(\mem~392_combout ),
	.datab(\mem~394_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~395_combout ),
	.cout());
defparam \mem~395 .lut_mask = 16'hAACC;
defparam \mem~395 .sum_lutc_input = "datac";

dffeas \internal_out_payload[22] (
	.clk(clk),
	.d(\mem~395_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[22]~q ),
	.prn(vcc));
defparam \internal_out_payload[22] .is_wysiwyg = "true";
defparam \internal_out_payload[22] .power_up = "low";

dffeas \mem~167 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~167_q ),
	.prn(vcc));
defparam \mem~167 .is_wysiwyg = "true";
defparam \mem~167 .power_up = "low";

dffeas \mem~199 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~199_q ),
	.prn(vcc));
defparam \mem~199 .is_wysiwyg = "true";
defparam \mem~199 .power_up = "low";

dffeas \mem~135 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~135_q ),
	.prn(vcc));
defparam \mem~135 .is_wysiwyg = "true";
defparam \mem~135 .power_up = "low";

cycloneive_lcell_comb \mem~396 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~199_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~135_q ),
	.cin(gnd),
	.combout(\mem~396_combout ),
	.cout());
defparam \mem~396 .lut_mask = 16'hFFDE;
defparam \mem~396 .sum_lutc_input = "datac";

dffeas \mem~231 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~231_q ),
	.prn(vcc));
defparam \mem~231 .is_wysiwyg = "true";
defparam \mem~231 .power_up = "low";

cycloneive_lcell_comb \mem~397 (
	.dataa(\mem~167_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~396_combout ),
	.datad(\mem~231_q ),
	.cin(gnd),
	.combout(\mem~397_combout ),
	.cout());
defparam \mem~397 .lut_mask = 16'hFFBE;
defparam \mem~397 .sum_lutc_input = "datac";

dffeas \mem~71 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~71_q ),
	.prn(vcc));
defparam \mem~71 .is_wysiwyg = "true";
defparam \mem~71 .power_up = "low";

dffeas \mem~39 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~39_q ),
	.prn(vcc));
defparam \mem~39 .is_wysiwyg = "true";
defparam \mem~39 .power_up = "low";

dffeas \mem~7 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~7_q ),
	.prn(vcc));
defparam \mem~7 .is_wysiwyg = "true";
defparam \mem~7 .power_up = "low";

cycloneive_lcell_comb \mem~398 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~39_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~7_q ),
	.cin(gnd),
	.combout(\mem~398_combout ),
	.cout());
defparam \mem~398 .lut_mask = 16'hFFDE;
defparam \mem~398 .sum_lutc_input = "datac";

dffeas \mem~103 (
	.clk(clk),
	.d(za_data_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~103_q ),
	.prn(vcc));
defparam \mem~103 .is_wysiwyg = "true";
defparam \mem~103 .power_up = "low";

cycloneive_lcell_comb \mem~399 (
	.dataa(\mem~71_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~398_combout ),
	.datad(\mem~103_q ),
	.cin(gnd),
	.combout(\mem~399_combout ),
	.cout());
defparam \mem~399 .lut_mask = 16'hFFBE;
defparam \mem~399 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~400 (
	.dataa(\mem~397_combout ),
	.datab(\mem~399_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~400_combout ),
	.cout());
defparam \mem~400 .lut_mask = 16'hAACC;
defparam \mem~400 .sum_lutc_input = "datac";

dffeas \internal_out_payload[7] (
	.clk(clk),
	.d(\mem~400_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[7]~q ),
	.prn(vcc));
defparam \internal_out_payload[7] .is_wysiwyg = "true";
defparam \internal_out_payload[7] .power_up = "low";

dffeas \mem~166 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~166_q ),
	.prn(vcc));
defparam \mem~166 .is_wysiwyg = "true";
defparam \mem~166 .power_up = "low";

dffeas \mem~198 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~198_q ),
	.prn(vcc));
defparam \mem~198 .is_wysiwyg = "true";
defparam \mem~198 .power_up = "low";

dffeas \mem~134 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~134_q ),
	.prn(vcc));
defparam \mem~134 .is_wysiwyg = "true";
defparam \mem~134 .power_up = "low";

cycloneive_lcell_comb \mem~401 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~198_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~134_q ),
	.cin(gnd),
	.combout(\mem~401_combout ),
	.cout());
defparam \mem~401 .lut_mask = 16'hFFDE;
defparam \mem~401 .sum_lutc_input = "datac";

dffeas \mem~230 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~230_q ),
	.prn(vcc));
defparam \mem~230 .is_wysiwyg = "true";
defparam \mem~230 .power_up = "low";

cycloneive_lcell_comb \mem~402 (
	.dataa(\mem~166_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~401_combout ),
	.datad(\mem~230_q ),
	.cin(gnd),
	.combout(\mem~402_combout ),
	.cout());
defparam \mem~402 .lut_mask = 16'hFFBE;
defparam \mem~402 .sum_lutc_input = "datac";

dffeas \mem~70 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~70_q ),
	.prn(vcc));
defparam \mem~70 .is_wysiwyg = "true";
defparam \mem~70 .power_up = "low";

dffeas \mem~38 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~38_q ),
	.prn(vcc));
defparam \mem~38 .is_wysiwyg = "true";
defparam \mem~38 .power_up = "low";

dffeas \mem~6 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~6_q ),
	.prn(vcc));
defparam \mem~6 .is_wysiwyg = "true";
defparam \mem~6 .power_up = "low";

cycloneive_lcell_comb \mem~403 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~38_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~6_q ),
	.cin(gnd),
	.combout(\mem~403_combout ),
	.cout());
defparam \mem~403 .lut_mask = 16'hFFDE;
defparam \mem~403 .sum_lutc_input = "datac";

dffeas \mem~102 (
	.clk(clk),
	.d(za_data_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~102_q ),
	.prn(vcc));
defparam \mem~102 .is_wysiwyg = "true";
defparam \mem~102 .power_up = "low";

cycloneive_lcell_comb \mem~404 (
	.dataa(\mem~70_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~403_combout ),
	.datad(\mem~102_q ),
	.cin(gnd),
	.combout(\mem~404_combout ),
	.cout());
defparam \mem~404 .lut_mask = 16'hFFBE;
defparam \mem~404 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~405 (
	.dataa(\mem~402_combout ),
	.datab(\mem~404_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~405_combout ),
	.cout());
defparam \mem~405 .lut_mask = 16'hAACC;
defparam \mem~405 .sum_lutc_input = "datac";

dffeas \internal_out_payload[6] (
	.clk(clk),
	.d(\mem~405_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[6]~q ),
	.prn(vcc));
defparam \internal_out_payload[6] .is_wysiwyg = "true";
defparam \internal_out_payload[6] .power_up = "low";

dffeas \mem~180 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~180_q ),
	.prn(vcc));
defparam \mem~180 .is_wysiwyg = "true";
defparam \mem~180 .power_up = "low";

dffeas \mem~212 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~212_q ),
	.prn(vcc));
defparam \mem~212 .is_wysiwyg = "true";
defparam \mem~212 .power_up = "low";

dffeas \mem~148 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~148_q ),
	.prn(vcc));
defparam \mem~148 .is_wysiwyg = "true";
defparam \mem~148 .power_up = "low";

cycloneive_lcell_comb \mem~406 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~212_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~148_q ),
	.cin(gnd),
	.combout(\mem~406_combout ),
	.cout());
defparam \mem~406 .lut_mask = 16'hFFDE;
defparam \mem~406 .sum_lutc_input = "datac";

dffeas \mem~244 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~244_q ),
	.prn(vcc));
defparam \mem~244 .is_wysiwyg = "true";
defparam \mem~244 .power_up = "low";

cycloneive_lcell_comb \mem~407 (
	.dataa(\mem~180_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~406_combout ),
	.datad(\mem~244_q ),
	.cin(gnd),
	.combout(\mem~407_combout ),
	.cout());
defparam \mem~407 .lut_mask = 16'hFFBE;
defparam \mem~407 .sum_lutc_input = "datac";

dffeas \mem~84 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~84_q ),
	.prn(vcc));
defparam \mem~84 .is_wysiwyg = "true";
defparam \mem~84 .power_up = "low";

dffeas \mem~52 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~52_q ),
	.prn(vcc));
defparam \mem~52 .is_wysiwyg = "true";
defparam \mem~52 .power_up = "low";

dffeas \mem~20 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~20_q ),
	.prn(vcc));
defparam \mem~20 .is_wysiwyg = "true";
defparam \mem~20 .power_up = "low";

cycloneive_lcell_comb \mem~408 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~52_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~20_q ),
	.cin(gnd),
	.combout(\mem~408_combout ),
	.cout());
defparam \mem~408 .lut_mask = 16'hFFDE;
defparam \mem~408 .sum_lutc_input = "datac";

dffeas \mem~116 (
	.clk(clk),
	.d(za_data_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~116_q ),
	.prn(vcc));
defparam \mem~116 .is_wysiwyg = "true";
defparam \mem~116 .power_up = "low";

cycloneive_lcell_comb \mem~409 (
	.dataa(\mem~84_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~408_combout ),
	.datad(\mem~116_q ),
	.cin(gnd),
	.combout(\mem~409_combout ),
	.cout());
defparam \mem~409 .lut_mask = 16'hFFBE;
defparam \mem~409 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~410 (
	.dataa(\mem~407_combout ),
	.datab(\mem~409_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~410_combout ),
	.cout());
defparam \mem~410 .lut_mask = 16'hAACC;
defparam \mem~410 .sum_lutc_input = "datac";

dffeas \internal_out_payload[20] (
	.clk(clk),
	.d(\mem~410_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[20]~q ),
	.prn(vcc));
defparam \internal_out_payload[20] .is_wysiwyg = "true";
defparam \internal_out_payload[20] .power_up = "low";

dffeas \mem~179 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~416_combout ),
	.q(\mem~179_q ),
	.prn(vcc));
defparam \mem~179 .is_wysiwyg = "true";
defparam \mem~179 .power_up = "low";

dffeas \mem~211 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~417_combout ),
	.q(\mem~211_q ),
	.prn(vcc));
defparam \mem~211 .is_wysiwyg = "true";
defparam \mem~211 .power_up = "low";

dffeas \mem~147 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~418_combout ),
	.q(\mem~147_q ),
	.prn(vcc));
defparam \mem~147 .is_wysiwyg = "true";
defparam \mem~147 .power_up = "low";

cycloneive_lcell_comb \mem~411 (
	.dataa(\mem_rd_ptr[0]~1_combout ),
	.datab(\mem~211_q ),
	.datac(\mem_rd_ptr[1]~0_combout ),
	.datad(\mem~147_q ),
	.cin(gnd),
	.combout(\mem~411_combout ),
	.cout());
defparam \mem~411 .lut_mask = 16'hFFDE;
defparam \mem~411 .sum_lutc_input = "datac";

dffeas \mem~243 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~419_combout ),
	.q(\mem~243_q ),
	.prn(vcc));
defparam \mem~243 .is_wysiwyg = "true";
defparam \mem~243 .power_up = "low";

cycloneive_lcell_comb \mem~412 (
	.dataa(\mem~179_q ),
	.datab(\mem_rd_ptr[0]~1_combout ),
	.datac(\mem~411_combout ),
	.datad(\mem~243_q ),
	.cin(gnd),
	.combout(\mem~412_combout ),
	.cout());
defparam \mem~412 .lut_mask = 16'hFFBE;
defparam \mem~412 .sum_lutc_input = "datac";

dffeas \mem~83 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~420_combout ),
	.q(\mem~83_q ),
	.prn(vcc));
defparam \mem~83 .is_wysiwyg = "true";
defparam \mem~83 .power_up = "low";

dffeas \mem~51 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~421_combout ),
	.q(\mem~51_q ),
	.prn(vcc));
defparam \mem~51 .is_wysiwyg = "true";
defparam \mem~51 .power_up = "low";

dffeas \mem~19 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~422_combout ),
	.q(\mem~19_q ),
	.prn(vcc));
defparam \mem~19 .is_wysiwyg = "true";
defparam \mem~19 .power_up = "low";

cycloneive_lcell_comb \mem~413 (
	.dataa(\mem_rd_ptr[1]~0_combout ),
	.datab(\mem~51_q ),
	.datac(\mem_rd_ptr[0]~1_combout ),
	.datad(\mem~19_q ),
	.cin(gnd),
	.combout(\mem~413_combout ),
	.cout());
defparam \mem~413 .lut_mask = 16'hFFDE;
defparam \mem~413 .sum_lutc_input = "datac";

dffeas \mem~115 (
	.clk(clk),
	.d(za_data_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem~423_combout ),
	.q(\mem~115_q ),
	.prn(vcc));
defparam \mem~115 .is_wysiwyg = "true";
defparam \mem~115 .power_up = "low";

cycloneive_lcell_comb \mem~414 (
	.dataa(\mem~83_q ),
	.datab(\mem_rd_ptr[1]~0_combout ),
	.datac(\mem~413_combout ),
	.datad(\mem~115_q ),
	.cin(gnd),
	.combout(\mem~414_combout ),
	.cout());
defparam \mem~414 .lut_mask = 16'hFFBE;
defparam \mem~414 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~415 (
	.dataa(\mem~412_combout ),
	.datab(\mem~414_combout ),
	.datac(gnd),
	.datad(\mem_rd_ptr[2]~2_combout ),
	.cin(gnd),
	.combout(\mem~415_combout ),
	.cout());
defparam \mem~415 .lut_mask = 16'hAACC;
defparam \mem~415 .sum_lutc_input = "datac";

dffeas \internal_out_payload[19] (
	.clk(clk),
	.d(\mem~415_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_payload[19]~q ),
	.prn(vcc));
defparam \internal_out_payload[19] .is_wysiwyg = "true";
defparam \internal_out_payload[19] .power_up = "low";

endmodule

module final_project_soc_altera_avalon_sc_fifo_10 (
	clk,
	reset,
	mem_used_7,
	last_cycle,
	saved_grant_0,
	saved_grant_1,
	WideOr1,
	out_data_buffer_67,
	src_data_68,
	nonposted_write_endofpacket,
	mem_used_0,
	mem_107_0,
	out_valid,
	mem_86_0,
	mem_68_0,
	WideOr0,
	mem_67_0,
	out_data_buffer_86)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
output 	mem_used_7;
input 	last_cycle;
input 	saved_grant_0;
input 	saved_grant_1;
input 	WideOr1;
input 	out_data_buffer_67;
input 	src_data_68;
input 	nonposted_write_endofpacket;
output 	mem_used_0;
output 	mem_107_0;
input 	out_valid;
output 	mem_86_0;
output 	mem_68_0;
input 	WideOr0;
output 	mem_67_0;
input 	out_data_buffer_86;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used~6_combout ;
wire \read~0_combout ;
wire \mem_used[6]~2_combout ;
wire \mem_used[1]~q ;
wire \mem_used~8_combout ;
wire \mem_used[2]~q ;
wire \mem_used~9_combout ;
wire \mem_used[3]~q ;
wire \mem_used~7_combout ;
wire \mem_used[4]~q ;
wire \mem_used~5_combout ;
wire \mem_used[5]~q ;
wire \mem_used~1_combout ;
wire \mem_used[6]~q ;
wire \mem_used[7]~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem[7][107]~q ;
wire \mem~24_combout ;
wire \always6~0_combout ;
wire \mem[6][107]~q ;
wire \mem~20_combout ;
wire \always5~0_combout ;
wire \mem[5][107]~q ;
wire \mem~16_combout ;
wire \always4~0_combout ;
wire \mem[4][107]~q ;
wire \mem~12_combout ;
wire \always3~0_combout ;
wire \mem[3][107]~q ;
wire \mem~8_combout ;
wire \always2~0_combout ;
wire \mem[2][107]~q ;
wire \mem~4_combout ;
wire \always1~0_combout ;
wire \mem[1][107]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[7][86]~q ;
wire \mem~25_combout ;
wire \mem[6][86]~q ;
wire \mem~21_combout ;
wire \mem[5][86]~q ;
wire \mem~17_combout ;
wire \mem[4][86]~q ;
wire \mem~13_combout ;
wire \mem[3][86]~q ;
wire \mem~9_combout ;
wire \mem[2][86]~q ;
wire \mem~5_combout ;
wire \mem[1][86]~q ;
wire \mem~1_combout ;
wire \mem[7][68]~q ;
wire \mem~26_combout ;
wire \mem[6][68]~q ;
wire \mem~22_combout ;
wire \mem[5][68]~q ;
wire \mem~18_combout ;
wire \mem[4][68]~q ;
wire \mem~14_combout ;
wire \mem[3][68]~q ;
wire \mem~10_combout ;
wire \mem[2][68]~q ;
wire \mem~6_combout ;
wire \mem[1][68]~q ;
wire \mem~2_combout ;
wire \mem[7][67]~q ;
wire \mem~27_combout ;
wire \mem[6][67]~q ;
wire \mem~23_combout ;
wire \mem[5][67]~q ;
wire \mem~19_combout ;
wire \mem[4][67]~q ;
wire \mem~15_combout ;
wire \mem[3][67]~q ;
wire \mem~11_combout ;
wire \mem[2][67]~q ;
wire \mem~7_combout ;
wire \mem[1][67]~q ;
wire \mem~3_combout ;


dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used[7]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_7),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(last_cycle),
	.datab(nonposted_write_endofpacket),
	.datac(WideOr1),
	.datad(src_data_68),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFFFE;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used~6 (
	.dataa(mem_used_0),
	.datab(\mem_used[2]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~6_combout ),
	.cout());
defparam \mem_used~6 .lut_mask = 16'hAACC;
defparam \mem_used~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(mem_used_0),
	.datab(mem_107_0),
	.datac(out_valid),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hFEFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[6]~2 (
	.dataa(\write~0_combout ),
	.datab(\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[6]~2_combout ),
	.cout());
defparam \mem_used[6]~2 .lut_mask = 16'h6666;
defparam \mem_used[6]~2 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used~8 (
	.dataa(\mem_used[1]~q ),
	.datab(\mem_used[3]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~8_combout ),
	.cout());
defparam \mem_used~8 .lut_mask = 16'hAACC;
defparam \mem_used~8 .sum_lutc_input = "datac";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cycloneive_lcell_comb \mem_used~9 (
	.dataa(\mem_used[2]~q ),
	.datab(\mem_used[4]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~9_combout ),
	.cout());
defparam \mem_used~9 .lut_mask = 16'hAACC;
defparam \mem_used~9 .sum_lutc_input = "datac";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cycloneive_lcell_comb \mem_used~7 (
	.dataa(\mem_used[3]~q ),
	.datab(\mem_used[5]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~7_combout ),
	.cout());
defparam \mem_used~7 .lut_mask = 16'hAACC;
defparam \mem_used~7 .sum_lutc_input = "datac";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cycloneive_lcell_comb \mem_used~5 (
	.dataa(\mem_used[4]~q ),
	.datab(\mem_used[6]~q ),
	.datac(gnd),
	.datad(\write~0_combout ),
	.cin(gnd),
	.combout(\mem_used~5_combout ),
	.cout());
defparam \mem_used~5 .lut_mask = 16'hAACC;
defparam \mem_used~5 .sum_lutc_input = "datac";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cycloneive_lcell_comb \mem_used~1 (
	.dataa(mem_used_7),
	.datab(\write~0_combout ),
	.datac(\mem_used[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used~1_combout ),
	.cout());
defparam \mem_used~1 .lut_mask = 16'hFEFE;
defparam \mem_used~1 .sum_lutc_input = "datac";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~2_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cycloneive_lcell_comb \mem_used[7]~0 (
	.dataa(mem_used_7),
	.datab(\write~0_combout ),
	.datac(\mem_used[6]~q ),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[7]~0_combout ),
	.cout());
defparam \mem_used[7]~0 .lut_mask = 16'hFBFE;
defparam \mem_used[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[1]~q ),
	.datab(gnd),
	.datac(mem_107_0),
	.datad(out_valid),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hAFFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\write~0_combout ),
	.datab(mem_used_0),
	.datac(WideOr0),
	.datad(\mem_used[0]~3_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem[7][107] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][107]~q ),
	.prn(vcc));
defparam \mem[7][107] .is_wysiwyg = "true";
defparam \mem[7][107] .power_up = "low";

cycloneive_lcell_comb \mem~24 (
	.dataa(\mem[7][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~24_combout ),
	.cout());
defparam \mem~24 .lut_mask = 16'hAACC;
defparam \mem~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always6~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\always6~0_combout ),
	.cout());
defparam \always6~0 .lut_mask = 16'hAAFF;
defparam \always6~0 .sum_lutc_input = "datac";

dffeas \mem[6][107] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][107]~q ),
	.prn(vcc));
defparam \mem[6][107] .is_wysiwyg = "true";
defparam \mem[6][107] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[6][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'hAAFF;
defparam \always5~0 .sum_lutc_input = "datac";

dffeas \mem[5][107] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][107]~q ),
	.prn(vcc));
defparam \mem[5][107] .is_wysiwyg = "true";
defparam \mem[5][107] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[5][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAACC;
defparam \mem~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hAAFF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas \mem[4][107] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][107]~q ),
	.prn(vcc));
defparam \mem[4][107] .is_wysiwyg = "true";
defparam \mem[4][107] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[4][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always3~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hAAFF;
defparam \always3~0 .sum_lutc_input = "datac";

dffeas \mem[3][107] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][107]~q ),
	.prn(vcc));
defparam \mem[3][107] .is_wysiwyg = "true";
defparam \mem[3][107] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[3][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hAACC;
defparam \mem~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

dffeas \mem[2][107] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][107]~q ),
	.prn(vcc));
defparam \mem[2][107] .is_wysiwyg = "true";
defparam \mem[2][107] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[2][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(\read~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hAAFF;
defparam \always1~0 .sum_lutc_input = "datac";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][107]~q ),
	.datab(nonposted_write_endofpacket),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(mem_107_0),
	.datab(out_valid),
	.datac(WideOr0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hEFFF;
defparam \always0~0 .sum_lutc_input = "datac";

dffeas \mem[7][86] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][86]~q ),
	.prn(vcc));
defparam \mem[7][86] .is_wysiwyg = "true";
defparam \mem[7][86] .power_up = "low";

cycloneive_lcell_comb \mem~25 (
	.dataa(\mem[7][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~25_combout ),
	.cout());
defparam \mem~25 .lut_mask = 16'hFAFC;
defparam \mem~25 .sum_lutc_input = "datac";

dffeas \mem[6][86] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][86]~q ),
	.prn(vcc));
defparam \mem[6][86] .is_wysiwyg = "true";
defparam \mem[6][86] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[6][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hFAFC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[5][86] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][86]~q ),
	.prn(vcc));
defparam \mem[5][86] .is_wysiwyg = "true";
defparam \mem[5][86] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[5][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hFAFC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[4][86] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][86]~q ),
	.prn(vcc));
defparam \mem[4][86] .is_wysiwyg = "true";
defparam \mem[4][86] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[4][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hFAFC;
defparam \mem~13 .sum_lutc_input = "datac";

dffeas \mem[3][86] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][86]~q ),
	.prn(vcc));
defparam \mem[3][86] .is_wysiwyg = "true";
defparam \mem[3][86] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[3][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hFAFC;
defparam \mem~9 .sum_lutc_input = "datac";

dffeas \mem[2][86] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][86]~q ),
	.prn(vcc));
defparam \mem[2][86] .is_wysiwyg = "true";
defparam \mem[2][86] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[2][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hFAFC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(out_data_buffer_86),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hFAFC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[7][68] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][68]~q ),
	.prn(vcc));
defparam \mem[7][68] .is_wysiwyg = "true";
defparam \mem[7][68] .power_up = "low";

cycloneive_lcell_comb \mem~26 (
	.dataa(\mem[7][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~26_combout ),
	.cout());
defparam \mem~26 .lut_mask = 16'hAACC;
defparam \mem~26 .sum_lutc_input = "datac";

dffeas \mem[6][68] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][68]~q ),
	.prn(vcc));
defparam \mem[6][68] .is_wysiwyg = "true";
defparam \mem[6][68] .power_up = "low";

cycloneive_lcell_comb \mem~22 (
	.dataa(\mem[6][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~22_combout ),
	.cout());
defparam \mem~22 .lut_mask = 16'hAACC;
defparam \mem~22 .sum_lutc_input = "datac";

dffeas \mem[5][68] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][68]~q ),
	.prn(vcc));
defparam \mem[5][68] .is_wysiwyg = "true";
defparam \mem[5][68] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[5][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

dffeas \mem[4][68] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][68]~q ),
	.prn(vcc));
defparam \mem[4][68] .is_wysiwyg = "true";
defparam \mem[4][68] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[4][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[3][68] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][68]~q ),
	.prn(vcc));
defparam \mem[3][68] .is_wysiwyg = "true";
defparam \mem[3][68] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[3][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hAACC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[2][68] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][68]~q ),
	.prn(vcc));
defparam \mem[2][68] .is_wysiwyg = "true";
defparam \mem[2][68] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[2][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[7][67] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][67]~q ),
	.prn(vcc));
defparam \mem[7][67] .is_wysiwyg = "true";
defparam \mem[7][67] .power_up = "low";

cycloneive_lcell_comb \mem~27 (
	.dataa(\mem[7][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(\mem~27_combout ),
	.cout());
defparam \mem~27 .lut_mask = 16'hFAFC;
defparam \mem~27 .sum_lutc_input = "datac";

dffeas \mem[6][67] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][67]~q ),
	.prn(vcc));
defparam \mem[6][67] .is_wysiwyg = "true";
defparam \mem[6][67] .power_up = "low";

cycloneive_lcell_comb \mem~23 (
	.dataa(\mem[6][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~23_combout ),
	.cout());
defparam \mem~23 .lut_mask = 16'hFAFC;
defparam \mem~23 .sum_lutc_input = "datac";

dffeas \mem[5][67] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][67]~q ),
	.prn(vcc));
defparam \mem[5][67] .is_wysiwyg = "true";
defparam \mem[5][67] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[5][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hFAFC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[4][67] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][67]~q ),
	.prn(vcc));
defparam \mem[4][67] .is_wysiwyg = "true";
defparam \mem[4][67] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[4][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hFAFC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[3][67] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][67]~q ),
	.prn(vcc));
defparam \mem[3][67] .is_wysiwyg = "true";
defparam \mem[3][67] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[3][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hFAFC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[2][67] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][67]~q ),
	.prn(vcc));
defparam \mem[2][67] .is_wysiwyg = "true";
defparam \mem[2][67] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[2][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hFAFC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][67]~q ),
	.datab(saved_grant_0),
	.datac(out_data_buffer_67),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hFAFC;
defparam \mem~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_sc_fifo_11 (
	uav_write,
	reset,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	mem_67_0,
	saved_grant_0,
	mem_used_1,
	saved_grant_1,
	WideOr1,
	cp_ready,
	src_data_68,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	uav_write;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_86_0;
output 	mem_68_0;
output 	mem_67_0;
input 	saved_grant_0;
output 	mem_used_1;
input 	saved_grant_1;
input 	WideOr1;
input 	cp_ready;
input 	src_data_68;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][86]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~1_combout ;
wire \mem[1][67]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem[0][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_86_0),
	.prn(vcc));
defparam \mem[0][86] .is_wysiwyg = "true";
defparam \mem[0][86] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[1][86] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][86]~q ),
	.prn(vcc));
defparam \mem[1][86] .is_wysiwyg = "true";
defparam \mem[1][86] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][86]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~2_combout ),
	.datab(WideOr1),
	.datac(src_data_68),
	.datad(cp_ready),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][68]~q ),
	.datab(src_data_68),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][67]~q ),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hFAFC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hACFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser (
	W_alu_result_4,
	W_alu_result_2,
	W_alu_result_3,
	clk_0,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	cp_valid,
	uav_write,
	d_writedata_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	uav_read,
	Equal3,
	take_in_data,
	saved_grant_0,
	out_data_buffer_3,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_buffer_67,
	out_data_buffer_31,
	out_data_buffer_107,
	mem_used_0,
	out_data_buffer_66,
	out_data_buffer_68,
	out_data_buffer_30,
	d_writedata_21,
	d_writedata_18,
	d_writedata_23,
	d_writedata_22,
	d_writedata_20,
	d_writedata_19,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_16,
	out_data_buffer_15,
	out_data_buffer_14,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_11,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_5,
	out_data_buffer_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	clk_0;
input 	d_writedata_31;
input 	d_writedata_30;
input 	d_writedata_29;
input 	d_writedata_28;
input 	d_writedata_27;
input 	d_writedata_26;
input 	d_writedata_25;
input 	d_writedata_24;
input 	cp_valid;
input 	uav_write;
input 	d_writedata_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	uav_read;
input 	Equal3;
output 	take_in_data;
input 	saved_grant_0;
output 	out_data_buffer_3;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
output 	out_data_buffer_67;
output 	out_data_buffer_31;
output 	out_data_buffer_107;
input 	mem_used_0;
output 	out_data_buffer_66;
output 	out_data_buffer_68;
output 	out_data_buffer_30;
input 	d_writedata_21;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_22;
input 	d_writedata_20;
input 	d_writedata_19;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_16;
output 	out_data_buffer_15;
output 	out_data_buffer_14;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_11;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_5;
output 	out_data_buffer_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_7 clock_xer(
	.W_alu_result_4(W_alu_result_4),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,uav_write,uav_write,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
W_alu_result_3,W_alu_result_2,gnd,gnd,gnd,gnd,gnd,gnd,d_writedata_31,d_writedata_30,d_writedata_29,d_writedata_28,d_writedata_27,d_writedata_26,d_writedata_25,d_writedata_24,d_writedata_23,d_writedata_22,d_writedata_21,d_writedata_20,d_writedata_19,d_writedata_18,d_writedata_17,
d_writedata_16,d_writedata_15,d_writedata_14,d_writedata_13,d_writedata_12,d_writedata_11,d_writedata_10,d_writedata_9,d_writedata_8,d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.clk_0(clk_0),
	.cp_valid(cp_valid),
	.in_reset(r_sync_rst),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.Equal3(Equal3),
	.take_in_data1(take_in_data),
	.saved_grant_0(saved_grant_0),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_107(out_data_buffer_107),
	.mem_used_0(mem_used_0),
	.out_data_buffer_66(out_data_buffer_66),
	.out_data_buffer_68(out_data_buffer_68),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_4(out_data_buffer_4),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_1 (
	wire_pll7_clk_0,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_11,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	cp_valid,
	uav_write,
	d_writedata_0,
	d_byteenable_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	altera_reset_synchronizer_int_chain_out,
	uav_read,
	in_ready,
	WideOr0,
	last_cycle,
	saved_grant_0,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_buffer_67,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	out_data_buffer_107,
	out_data_buffer_66,
	d_byteenable_2,
	WideOr01,
	d_byteenable_1,
	d_byteenable_3,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_18,
	out_data_buffer_19,
	out_data_buffer_20,
	out_data_buffer_21,
	out_data_buffer_22,
	out_data_buffer_23,
	out_data_buffer_24,
	out_data_buffer_25,
	out_data_buffer_26,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_29,
	out_data_buffer_30,
	out_data_buffer_31,
	d_writedata_21,
	d_writedata_18,
	d_writedata_23,
	d_writedata_22,
	d_writedata_20,
	d_writedata_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_24;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_12;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_11;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_31;
input 	d_writedata_30;
input 	d_writedata_29;
input 	d_writedata_28;
input 	d_writedata_27;
input 	d_writedata_26;
input 	d_writedata_25;
input 	d_writedata_24;
input 	cp_valid;
input 	uav_write;
input 	d_writedata_0;
input 	d_byteenable_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	altera_reset_synchronizer_int_chain_out;
input 	uav_read;
output 	in_ready;
input 	WideOr0;
input 	last_cycle;
input 	saved_grant_0;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
output 	out_data_buffer_67;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
output 	out_data_buffer_107;
output 	out_data_buffer_66;
input 	d_byteenable_2;
input 	WideOr01;
input 	d_byteenable_1;
input 	d_byteenable_3;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_18;
output 	out_data_buffer_19;
output 	out_data_buffer_20;
output 	out_data_buffer_21;
output 	out_data_buffer_22;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_29;
output 	out_data_buffer_30;
output 	out_data_buffer_31;
input 	d_writedata_21;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_22;
input 	d_writedata_20;
input 	d_writedata_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,uav_read,uav_write,uav_write,gnd,gnd,gnd,W_alu_result_26,W_alu_result_25,W_alu_result_24,W_alu_result_23,
W_alu_result_22,W_alu_result_21,W_alu_result_20,W_alu_result_19,W_alu_result_18,W_alu_result_17,W_alu_result_16,W_alu_result_15,W_alu_result_14,W_alu_result_13,W_alu_result_12,W_alu_result_11,W_alu_result_10,W_alu_result_9,W_alu_result_8,W_alu_result_7,W_alu_result_6,
W_alu_result_5,W_alu_result_4,W_alu_result_3,W_alu_result_2,gnd,gnd,d_byteenable_3,d_byteenable_2,d_byteenable_1,d_byteenable_0,d_writedata_31,d_writedata_30,d_writedata_29,d_writedata_28,d_writedata_27,d_writedata_26,d_writedata_25,d_writedata_24,d_writedata_23,
d_writedata_22,d_writedata_21,d_writedata_20,d_writedata_19,d_writedata_18,d_writedata_17,d_writedata_16,d_writedata_15,d_writedata_14,d_writedata_13,d_writedata_12,d_writedata_11,d_writedata_10,d_writedata_9,d_writedata_8,d_writedata_7,d_writedata_6,d_writedata_5,
d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.cp_valid(cp_valid),
	.in_reset(r_sync_rst),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.in_ready(in_ready),
	.WideOr0(WideOr0),
	.last_cycle(last_cycle),
	.saved_grant_0(saved_grant_0),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_68(out_data_buffer_68),
	.out_data_buffer_48(out_data_buffer_48),
	.out_data_buffer_62(out_data_buffer_62),
	.out_data_buffer_49(out_data_buffer_49),
	.out_data_buffer_51(out_data_buffer_51),
	.out_data_buffer_50(out_data_buffer_50),
	.out_data_buffer_53(out_data_buffer_53),
	.out_data_buffer_52(out_data_buffer_52),
	.out_data_buffer_55(out_data_buffer_55),
	.out_data_buffer_54(out_data_buffer_54),
	.out_data_buffer_57(out_data_buffer_57),
	.out_data_buffer_56(out_data_buffer_56),
	.out_data_buffer_59(out_data_buffer_59),
	.out_data_buffer_58(out_data_buffer_58),
	.out_data_buffer_61(out_data_buffer_61),
	.out_data_buffer_60(out_data_buffer_60),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_buffer_40(out_data_buffer_40),
	.out_data_buffer_41(out_data_buffer_41),
	.out_data_buffer_42(out_data_buffer_42),
	.out_data_buffer_43(out_data_buffer_43),
	.out_data_buffer_44(out_data_buffer_44),
	.out_data_buffer_45(out_data_buffer_45),
	.out_data_buffer_46(out_data_buffer_46),
	.out_data_buffer_47(out_data_buffer_47),
	.out_data_buffer_32(out_data_buffer_32),
	.out_data_buffer_33(out_data_buffer_33),
	.out_data_buffer_34(out_data_buffer_34),
	.out_data_buffer_35(out_data_buffer_35),
	.out_data_buffer_107(out_data_buffer_107),
	.out_data_buffer_66(out_data_buffer_66),
	.WideOr01(WideOr01),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_31(out_data_buffer_31),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser (
	wire_pll7_clk_0,
	in_data,
	cp_valid,
	in_reset,
	out_reset,
	in_ready,
	WideOr0,
	last_cycle,
	saved_grant_0,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	out_data_buffer_67,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	out_data_buffer_107,
	out_data_buffer_66,
	WideOr01,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_18,
	out_data_buffer_19,
	out_data_buffer_20,
	out_data_buffer_21,
	out_data_buffer_22,
	out_data_buffer_23,
	out_data_buffer_24,
	out_data_buffer_25,
	out_data_buffer_26,
	out_data_buffer_27,
	out_data_buffer_28,
	out_data_buffer_29,
	out_data_buffer_30,
	out_data_buffer_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	[118:0] in_data;
input 	cp_valid;
input 	in_reset;
input 	out_reset;
output 	in_ready;
input 	WideOr0;
input 	last_cycle;
input 	saved_grant_0;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
output 	out_data_buffer_67;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
output 	out_data_buffer_107;
output 	out_data_buffer_66;
input 	WideOr01;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_18;
output 	out_data_buffer_19;
output 	out_data_buffer_20;
output 	out_data_buffer_21;
output 	out_data_buffer_22;
output 	out_data_buffer_23;
output 	out_data_buffer_24;
output 	out_data_buffer_25;
output 	out_data_buffer_26;
output 	out_data_buffer_27;
output 	out_data_buffer_28;
output 	out_data_buffer_29;
output 	out_data_buffer_30;
output 	out_data_buffer_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_toggle~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \take_in_data~0_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_buffer[68]~q ;
wire \in_data_buffer[48]~q ;
wire \in_data_buffer[62]~q ;
wire \in_data_buffer[49]~q ;
wire \in_data_buffer[51]~q ;
wire \in_data_buffer[50]~q ;
wire \in_data_buffer[53]~q ;
wire \in_data_buffer[52]~q ;
wire \in_data_buffer[55]~q ;
wire \in_data_buffer[54]~q ;
wire \in_data_buffer[57]~q ;
wire \in_data_buffer[56]~q ;
wire \in_data_buffer[59]~q ;
wire \in_data_buffer[58]~q ;
wire \in_data_buffer[61]~q ;
wire \in_data_buffer[60]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[40]~q ;
wire \in_data_buffer[41]~q ;
wire \in_data_buffer[42]~q ;
wire \in_data_buffer[43]~q ;
wire \in_data_buffer[44]~q ;
wire \in_data_buffer[45]~q ;
wire \in_data_buffer[46]~q ;
wire \in_data_buffer[47]~q ;
wire \in_data_buffer[32]~q ;
wire \in_data_buffer[33]~q ;
wire \in_data_buffer[34]~q ;
wire \in_data_buffer[35]~q ;
wire \in_data_buffer[107]~q ;
wire \in_data_buffer[66]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[31]~q ;


final_project_soc_altera_std_synchronizer_2 out_to_in_synchronizer(
	.reset_n(in_reset),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ),
	.din(out_data_toggle_flopped1),
	.clk(clk_clk));

final_project_soc_altera_std_synchronizer_1 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.din(\in_data_toggle~q ),
	.dreg_0(dreg_0));

cycloneive_lcell_comb \in_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(in_ready),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h0FF0;
defparam \in_ready~0 .sum_lutc_input = "datac";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas \out_data_buffer[68] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[68]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_68),
	.prn(vcc));
defparam \out_data_buffer[68] .is_wysiwyg = "true";
defparam \out_data_buffer[68] .power_up = "low";

dffeas \out_data_buffer[48] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[48]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_48),
	.prn(vcc));
defparam \out_data_buffer[48] .is_wysiwyg = "true";
defparam \out_data_buffer[48] .power_up = "low";

dffeas \out_data_buffer[62] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[62]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_62),
	.prn(vcc));
defparam \out_data_buffer[62] .is_wysiwyg = "true";
defparam \out_data_buffer[62] .power_up = "low";

dffeas \out_data_buffer[49] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[49]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_49),
	.prn(vcc));
defparam \out_data_buffer[49] .is_wysiwyg = "true";
defparam \out_data_buffer[49] .power_up = "low";

dffeas \out_data_buffer[51] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[51]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_51),
	.prn(vcc));
defparam \out_data_buffer[51] .is_wysiwyg = "true";
defparam \out_data_buffer[51] .power_up = "low";

dffeas \out_data_buffer[50] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[50]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_50),
	.prn(vcc));
defparam \out_data_buffer[50] .is_wysiwyg = "true";
defparam \out_data_buffer[50] .power_up = "low";

dffeas \out_data_buffer[53] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[53]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_53),
	.prn(vcc));
defparam \out_data_buffer[53] .is_wysiwyg = "true";
defparam \out_data_buffer[53] .power_up = "low";

dffeas \out_data_buffer[52] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[52]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_52),
	.prn(vcc));
defparam \out_data_buffer[52] .is_wysiwyg = "true";
defparam \out_data_buffer[52] .power_up = "low";

dffeas \out_data_buffer[55] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[55]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_55),
	.prn(vcc));
defparam \out_data_buffer[55] .is_wysiwyg = "true";
defparam \out_data_buffer[55] .power_up = "low";

dffeas \out_data_buffer[54] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[54]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_54),
	.prn(vcc));
defparam \out_data_buffer[54] .is_wysiwyg = "true";
defparam \out_data_buffer[54] .power_up = "low";

dffeas \out_data_buffer[57] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[57]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_57),
	.prn(vcc));
defparam \out_data_buffer[57] .is_wysiwyg = "true";
defparam \out_data_buffer[57] .power_up = "low";

dffeas \out_data_buffer[56] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[56]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_56),
	.prn(vcc));
defparam \out_data_buffer[56] .is_wysiwyg = "true";
defparam \out_data_buffer[56] .power_up = "low";

dffeas \out_data_buffer[59] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[59]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_59),
	.prn(vcc));
defparam \out_data_buffer[59] .is_wysiwyg = "true";
defparam \out_data_buffer[59] .power_up = "low";

dffeas \out_data_buffer[58] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[58]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_58),
	.prn(vcc));
defparam \out_data_buffer[58] .is_wysiwyg = "true";
defparam \out_data_buffer[58] .power_up = "low";

dffeas \out_data_buffer[61] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[61]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_61),
	.prn(vcc));
defparam \out_data_buffer[61] .is_wysiwyg = "true";
defparam \out_data_buffer[61] .power_up = "low";

dffeas \out_data_buffer[60] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[60]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_60),
	.prn(vcc));
defparam \out_data_buffer[60] .is_wysiwyg = "true";
defparam \out_data_buffer[60] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas \out_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[40]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_40),
	.prn(vcc));
defparam \out_data_buffer[40] .is_wysiwyg = "true";
defparam \out_data_buffer[40] .power_up = "low";

dffeas \out_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[41]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_41),
	.prn(vcc));
defparam \out_data_buffer[41] .is_wysiwyg = "true";
defparam \out_data_buffer[41] .power_up = "low";

dffeas \out_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[42]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_42),
	.prn(vcc));
defparam \out_data_buffer[42] .is_wysiwyg = "true";
defparam \out_data_buffer[42] .power_up = "low";

dffeas \out_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[43]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_43),
	.prn(vcc));
defparam \out_data_buffer[43] .is_wysiwyg = "true";
defparam \out_data_buffer[43] .power_up = "low";

dffeas \out_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[44]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_44),
	.prn(vcc));
defparam \out_data_buffer[44] .is_wysiwyg = "true";
defparam \out_data_buffer[44] .power_up = "low";

dffeas \out_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[45]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_45),
	.prn(vcc));
defparam \out_data_buffer[45] .is_wysiwyg = "true";
defparam \out_data_buffer[45] .power_up = "low";

dffeas \out_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[46]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_46),
	.prn(vcc));
defparam \out_data_buffer[46] .is_wysiwyg = "true";
defparam \out_data_buffer[46] .power_up = "low";

dffeas \out_data_buffer[47] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[47]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_47),
	.prn(vcc));
defparam \out_data_buffer[47] .is_wysiwyg = "true";
defparam \out_data_buffer[47] .power_up = "low";

dffeas \out_data_buffer[32] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[32]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_32),
	.prn(vcc));
defparam \out_data_buffer[32] .is_wysiwyg = "true";
defparam \out_data_buffer[32] .power_up = "low";

dffeas \out_data_buffer[33] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[33]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_33),
	.prn(vcc));
defparam \out_data_buffer[33] .is_wysiwyg = "true";
defparam \out_data_buffer[33] .power_up = "low";

dffeas \out_data_buffer[34] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[34]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_34),
	.prn(vcc));
defparam \out_data_buffer[34] .is_wysiwyg = "true";
defparam \out_data_buffer[34] .power_up = "low";

dffeas \out_data_buffer[35] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[35]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_35),
	.prn(vcc));
defparam \out_data_buffer[35] .is_wysiwyg = "true";
defparam \out_data_buffer[35] .power_up = "low";

dffeas \out_data_buffer[107] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[107]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_107),
	.prn(vcc));
defparam \out_data_buffer[107] .is_wysiwyg = "true";
defparam \out_data_buffer[107] .power_up = "low";

dffeas \out_data_buffer[66] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(gnd),
	.datab(\in_data_toggle~q ),
	.datac(cp_valid),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hC33C;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(dreg_0),
	.datab(out_data_toggle_flopped1),
	.datac(last_cycle),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(cp_valid),
	.datab(WideOr01),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\take_in_data~0_combout ),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hEFFE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(clk_clk),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

dffeas \in_data_buffer[68] (
	.clk(clk_clk),
	.d(in_data[68]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[68]~q ),
	.prn(vcc));
defparam \in_data_buffer[68] .is_wysiwyg = "true";
defparam \in_data_buffer[68] .power_up = "low";

dffeas \in_data_buffer[48] (
	.clk(clk_clk),
	.d(in_data[48]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[48]~q ),
	.prn(vcc));
defparam \in_data_buffer[48] .is_wysiwyg = "true";
defparam \in_data_buffer[48] .power_up = "low";

dffeas \in_data_buffer[62] (
	.clk(clk_clk),
	.d(in_data[62]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[62]~q ),
	.prn(vcc));
defparam \in_data_buffer[62] .is_wysiwyg = "true";
defparam \in_data_buffer[62] .power_up = "low";

dffeas \in_data_buffer[49] (
	.clk(clk_clk),
	.d(in_data[49]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[49]~q ),
	.prn(vcc));
defparam \in_data_buffer[49] .is_wysiwyg = "true";
defparam \in_data_buffer[49] .power_up = "low";

dffeas \in_data_buffer[51] (
	.clk(clk_clk),
	.d(in_data[51]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[51]~q ),
	.prn(vcc));
defparam \in_data_buffer[51] .is_wysiwyg = "true";
defparam \in_data_buffer[51] .power_up = "low";

dffeas \in_data_buffer[50] (
	.clk(clk_clk),
	.d(in_data[50]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[50]~q ),
	.prn(vcc));
defparam \in_data_buffer[50] .is_wysiwyg = "true";
defparam \in_data_buffer[50] .power_up = "low";

dffeas \in_data_buffer[53] (
	.clk(clk_clk),
	.d(in_data[53]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[53]~q ),
	.prn(vcc));
defparam \in_data_buffer[53] .is_wysiwyg = "true";
defparam \in_data_buffer[53] .power_up = "low";

dffeas \in_data_buffer[52] (
	.clk(clk_clk),
	.d(in_data[52]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[52]~q ),
	.prn(vcc));
defparam \in_data_buffer[52] .is_wysiwyg = "true";
defparam \in_data_buffer[52] .power_up = "low";

dffeas \in_data_buffer[55] (
	.clk(clk_clk),
	.d(in_data[55]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[55]~q ),
	.prn(vcc));
defparam \in_data_buffer[55] .is_wysiwyg = "true";
defparam \in_data_buffer[55] .power_up = "low";

dffeas \in_data_buffer[54] (
	.clk(clk_clk),
	.d(in_data[54]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[54]~q ),
	.prn(vcc));
defparam \in_data_buffer[54] .is_wysiwyg = "true";
defparam \in_data_buffer[54] .power_up = "low";

dffeas \in_data_buffer[57] (
	.clk(clk_clk),
	.d(in_data[57]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[57]~q ),
	.prn(vcc));
defparam \in_data_buffer[57] .is_wysiwyg = "true";
defparam \in_data_buffer[57] .power_up = "low";

dffeas \in_data_buffer[56] (
	.clk(clk_clk),
	.d(in_data[56]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[56]~q ),
	.prn(vcc));
defparam \in_data_buffer[56] .is_wysiwyg = "true";
defparam \in_data_buffer[56] .power_up = "low";

dffeas \in_data_buffer[59] (
	.clk(clk_clk),
	.d(in_data[59]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[59]~q ),
	.prn(vcc));
defparam \in_data_buffer[59] .is_wysiwyg = "true";
defparam \in_data_buffer[59] .power_up = "low";

dffeas \in_data_buffer[58] (
	.clk(clk_clk),
	.d(in_data[58]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[58]~q ),
	.prn(vcc));
defparam \in_data_buffer[58] .is_wysiwyg = "true";
defparam \in_data_buffer[58] .power_up = "low";

dffeas \in_data_buffer[61] (
	.clk(clk_clk),
	.d(in_data[61]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[61]~q ),
	.prn(vcc));
defparam \in_data_buffer[61] .is_wysiwyg = "true";
defparam \in_data_buffer[61] .power_up = "low";

dffeas \in_data_buffer[60] (
	.clk(clk_clk),
	.d(in_data[60]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[60]~q ),
	.prn(vcc));
defparam \in_data_buffer[60] .is_wysiwyg = "true";
defparam \in_data_buffer[60] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(clk_clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(clk_clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[40] (
	.clk(clk_clk),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[40]~q ),
	.prn(vcc));
defparam \in_data_buffer[40] .is_wysiwyg = "true";
defparam \in_data_buffer[40] .power_up = "low";

dffeas \in_data_buffer[41] (
	.clk(clk_clk),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[41]~q ),
	.prn(vcc));
defparam \in_data_buffer[41] .is_wysiwyg = "true";
defparam \in_data_buffer[41] .power_up = "low";

dffeas \in_data_buffer[42] (
	.clk(clk_clk),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[42]~q ),
	.prn(vcc));
defparam \in_data_buffer[42] .is_wysiwyg = "true";
defparam \in_data_buffer[42] .power_up = "low";

dffeas \in_data_buffer[43] (
	.clk(clk_clk),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[43]~q ),
	.prn(vcc));
defparam \in_data_buffer[43] .is_wysiwyg = "true";
defparam \in_data_buffer[43] .power_up = "low";

dffeas \in_data_buffer[44] (
	.clk(clk_clk),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[44]~q ),
	.prn(vcc));
defparam \in_data_buffer[44] .is_wysiwyg = "true";
defparam \in_data_buffer[44] .power_up = "low";

dffeas \in_data_buffer[45] (
	.clk(clk_clk),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[45]~q ),
	.prn(vcc));
defparam \in_data_buffer[45] .is_wysiwyg = "true";
defparam \in_data_buffer[45] .power_up = "low";

dffeas \in_data_buffer[46] (
	.clk(clk_clk),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[46]~q ),
	.prn(vcc));
defparam \in_data_buffer[46] .is_wysiwyg = "true";
defparam \in_data_buffer[46] .power_up = "low";

dffeas \in_data_buffer[47] (
	.clk(clk_clk),
	.d(in_data[47]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[47]~q ),
	.prn(vcc));
defparam \in_data_buffer[47] .is_wysiwyg = "true";
defparam \in_data_buffer[47] .power_up = "low";

dffeas \in_data_buffer[32] (
	.clk(clk_clk),
	.d(in_data[32]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[32]~q ),
	.prn(vcc));
defparam \in_data_buffer[32] .is_wysiwyg = "true";
defparam \in_data_buffer[32] .power_up = "low";

dffeas \in_data_buffer[33] (
	.clk(clk_clk),
	.d(in_data[33]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[33]~q ),
	.prn(vcc));
defparam \in_data_buffer[33] .is_wysiwyg = "true";
defparam \in_data_buffer[33] .power_up = "low";

dffeas \in_data_buffer[34] (
	.clk(clk_clk),
	.d(in_data[34]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[34]~q ),
	.prn(vcc));
defparam \in_data_buffer[34] .is_wysiwyg = "true";
defparam \in_data_buffer[34] .power_up = "low";

dffeas \in_data_buffer[35] (
	.clk(clk_clk),
	.d(in_data[35]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[35]~q ),
	.prn(vcc));
defparam \in_data_buffer[35] .is_wysiwyg = "true";
defparam \in_data_buffer[35] .power_up = "low";

dffeas \in_data_buffer[107] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[107]~q ),
	.prn(vcc));
defparam \in_data_buffer[107] .is_wysiwyg = "true";
defparam \in_data_buffer[107] .power_up = "low";

dffeas \in_data_buffer[66] (
	.clk(clk_clk),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(clk_clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(clk_clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(clk_clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(clk_clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(clk_clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(clk_clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(clk_clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(clk_clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(clk_clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(clk_clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(clk_clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(clk_clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(clk_clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(clk_clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(clk_clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(clk_clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(clk_clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(clk_clk),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(clk_clk),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(clk_clk),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(clk_clk),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(clk_clk),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(clk_clk),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(clk_clk),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(clk_clk),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(clk_clk),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_1 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_2 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_2 (
	clk_0,
	i_read,
	read_accepted,
	F_pc_2,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	Equal2,
	take_in_data,
	saved_grant_1,
	out_data_buffer_38,
	out_data_buffer_39,
	out_valid,
	out_data_buffer_107,
	mem_used_0,
	out_data_buffer_68,
	out_data_buffer_86,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	i_read;
input 	read_accepted;
input 	F_pc_2;
input 	F_pc_0;
input 	F_pc_1;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal2;
output 	take_in_data;
input 	saved_grant_1;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_valid;
output 	out_data_buffer_107;
input 	mem_used_0;
output 	out_data_buffer_68;
output 	out_data_buffer_86;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_1 clock_xer(
	.clk_0(clk_0),
	.i_read(i_read),
	.read_accepted(read_accepted),
	.F_pc_2(F_pc_2),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,F_pc_1,F_pc_0,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.in_reset(r_sync_rst),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.Equal2(Equal2),
	.take_in_data1(take_in_data),
	.saved_grant_1(saved_grant_1),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_valid1(out_valid),
	.out_data_buffer_107(out_data_buffer_107),
	.mem_used_0(mem_used_0),
	.out_data_buffer_68(out_data_buffer_68),
	.out_data_buffer_86(out_data_buffer_86),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_1 (
	clk_0,
	i_read,
	read_accepted,
	F_pc_2,
	in_data,
	in_reset,
	out_reset,
	Equal2,
	take_in_data1,
	saved_grant_1,
	out_data_buffer_38,
	out_data_buffer_39,
	out_valid1,
	out_data_buffer_107,
	mem_used_0,
	out_data_buffer_68,
	out_data_buffer_86,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	i_read;
input 	read_accepted;
input 	F_pc_2;
input 	[118:0] in_data;
input 	in_reset;
input 	out_reset;
input 	Equal2;
output 	take_in_data1;
input 	saved_grant_1;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_valid1;
output 	out_data_buffer_107;
input 	mem_used_0;
output 	out_data_buffer_68;
output 	out_data_buffer_86;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_to_out_synchronizer|dreg[0]~q ;
wire \in_data_toggle~2_combout ;
wire \in_data_toggle~q ;
wire \take_in_data~combout ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \out_data_toggle_flopped~q ;
wire \in_data_buffer[107]~q ;
wire \in_data_buffer[68]~q ;
wire \in_data_buffer[86]~q ;


final_project_soc_altera_std_synchronizer_4 out_to_in_synchronizer(
	.reset_n(in_reset),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ),
	.din(\out_data_toggle_flopped~q ),
	.clk(clk_clk));

final_project_soc_altera_std_synchronizer_3 in_to_out_synchronizer(
	.clk(clk_0),
	.reset_n(out_reset),
	.din(\in_data_toggle~q ),
	.dreg_0(\in_to_out_synchronizer|dreg[0]~q ));

cycloneive_lcell_comb \take_in_data~2 (
	.dataa(Equal2),
	.datab(\in_data_toggle~q ),
	.datac(\out_to_in_synchronizer|dreg[0]~q ),
	.datad(F_pc_2),
	.cin(gnd),
	.combout(take_in_data1),
	.cout());
defparam \take_in_data~2 .lut_mask = 16'hBEFF;
defparam \take_in_data~2 .sum_lutc_input = "datac";

dffeas \out_data_buffer[38] (
	.clk(clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_data_toggle_flopped~q ),
	.datad(\in_to_out_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[107] (
	.clk(clk_0),
	.d(\in_data_buffer[107]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_107),
	.prn(vcc));
defparam \out_data_buffer[107] .is_wysiwyg = "true";
defparam \out_data_buffer[107] .power_up = "low";

dffeas \out_data_buffer[68] (
	.clk(clk_0),
	.d(\in_data_buffer[68]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_68),
	.prn(vcc));
defparam \out_data_buffer[68] .is_wysiwyg = "true";
defparam \out_data_buffer[68] .power_up = "low";

dffeas \out_data_buffer[86] (
	.clk(clk_0),
	.d(\in_data_buffer[86]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_86),
	.prn(vcc));
defparam \out_data_buffer[86] .is_wysiwyg = "true";
defparam \out_data_buffer[86] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(\in_data_toggle~q ),
	.datad(take_in_data1),
	.cin(gnd),
	.combout(\in_data_toggle~2_combout ),
	.cout());
defparam \in_data_toggle~2 .lut_mask = 16'h6996;
defparam \in_data_toggle~2 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~2_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb take_in_data(
	.dataa(i_read),
	.datab(read_accepted),
	.datac(take_in_data1),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hF7F7;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[38] (
	.clk(clk_clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(clk_clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(\in_to_out_synchronizer|dreg[0]~q ),
	.datab(\out_data_toggle_flopped~q ),
	.datac(saved_grant_1),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas out_data_toggle_flopped(
	.clk(clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_toggle_flopped~q ),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

dffeas \in_data_buffer[107] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[107]~q ),
	.prn(vcc));
defparam \in_data_buffer[107] .is_wysiwyg = "true";
defparam \in_data_buffer[107] .power_up = "low";

dffeas \in_data_buffer[68] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[68]~q ),
	.prn(vcc));
defparam \in_data_buffer[68] .is_wysiwyg = "true";
defparam \in_data_buffer[68] .power_up = "low";

dffeas \in_data_buffer[86] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[86]~q ),
	.prn(vcc));
defparam \in_data_buffer[86] .is_wysiwyg = "true";
defparam \in_data_buffer[86] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_3 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_4 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_3 (
	wire_pll7_clk_0,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_3,
	uav_read,
	F_pc_2,
	F_pc_4,
	F_pc_9,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	src_channel_5,
	in_ready,
	last_cycle,
	saved_grant_1,
	out_valid,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	out_data_buffer_107,
	out_data_buffer_86,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	F_pc_10;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_3;
input 	uav_read;
input 	F_pc_2;
input 	F_pc_4;
input 	F_pc_9;
input 	F_pc_0;
input 	F_pc_1;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
input 	src_channel_5;
output 	in_ready;
input 	last_cycle;
input 	saved_grant_1;
output 	out_valid;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
output 	out_data_buffer_107;
output 	out_data_buffer_86;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_2 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,F_pc_24,F_pc_23,F_pc_22,F_pc_21,F_pc_20,F_pc_19,F_pc_18,F_pc_17,F_pc_16,F_pc_15,F_pc_14,F_pc_13,
F_pc_12,F_pc_11,F_pc_10,F_pc_9,F_pc_8,F_pc_7,F_pc_6,F_pc_5,F_pc_4,F_pc_3,F_pc_2,F_pc_1,F_pc_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.uav_read(uav_read),
	.in_reset(r_sync_rst),
	.out_reset(altera_reset_synchronizer_int_chain_out),
	.src_channel_5(src_channel_5),
	.in_ready(in_ready),
	.last_cycle(last_cycle),
	.saved_grant_1(saved_grant_1),
	.out_valid1(out_valid),
	.out_data_buffer_68(out_data_buffer_68),
	.out_data_buffer_48(out_data_buffer_48),
	.out_data_buffer_62(out_data_buffer_62),
	.out_data_buffer_49(out_data_buffer_49),
	.out_data_buffer_51(out_data_buffer_51),
	.out_data_buffer_50(out_data_buffer_50),
	.out_data_buffer_53(out_data_buffer_53),
	.out_data_buffer_52(out_data_buffer_52),
	.out_data_buffer_55(out_data_buffer_55),
	.out_data_buffer_54(out_data_buffer_54),
	.out_data_buffer_57(out_data_buffer_57),
	.out_data_buffer_56(out_data_buffer_56),
	.out_data_buffer_59(out_data_buffer_59),
	.out_data_buffer_58(out_data_buffer_58),
	.out_data_buffer_61(out_data_buffer_61),
	.out_data_buffer_60(out_data_buffer_60),
	.out_data_buffer_38(out_data_buffer_38),
	.out_data_buffer_39(out_data_buffer_39),
	.out_data_buffer_40(out_data_buffer_40),
	.out_data_buffer_41(out_data_buffer_41),
	.out_data_buffer_42(out_data_buffer_42),
	.out_data_buffer_43(out_data_buffer_43),
	.out_data_buffer_44(out_data_buffer_44),
	.out_data_buffer_45(out_data_buffer_45),
	.out_data_buffer_46(out_data_buffer_46),
	.out_data_buffer_47(out_data_buffer_47),
	.out_data_buffer_32(out_data_buffer_32),
	.out_data_buffer_33(out_data_buffer_33),
	.out_data_buffer_34(out_data_buffer_34),
	.out_data_buffer_35(out_data_buffer_35),
	.out_data_buffer_107(out_data_buffer_107),
	.out_data_buffer_86(out_data_buffer_86),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_2 (
	wire_pll7_clk_0,
	in_data,
	uav_read,
	in_reset,
	out_reset,
	src_channel_5,
	in_ready,
	last_cycle,
	saved_grant_1,
	out_valid1,
	out_data_buffer_68,
	out_data_buffer_48,
	out_data_buffer_62,
	out_data_buffer_49,
	out_data_buffer_51,
	out_data_buffer_50,
	out_data_buffer_53,
	out_data_buffer_52,
	out_data_buffer_55,
	out_data_buffer_54,
	out_data_buffer_57,
	out_data_buffer_56,
	out_data_buffer_59,
	out_data_buffer_58,
	out_data_buffer_61,
	out_data_buffer_60,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_buffer_40,
	out_data_buffer_41,
	out_data_buffer_42,
	out_data_buffer_43,
	out_data_buffer_44,
	out_data_buffer_45,
	out_data_buffer_46,
	out_data_buffer_47,
	out_data_buffer_32,
	out_data_buffer_33,
	out_data_buffer_34,
	out_data_buffer_35,
	out_data_buffer_107,
	out_data_buffer_86,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	[118:0] in_data;
input 	uav_read;
input 	in_reset;
input 	out_reset;
input 	src_channel_5;
output 	in_ready;
input 	last_cycle;
input 	saved_grant_1;
output 	out_valid1;
output 	out_data_buffer_68;
output 	out_data_buffer_48;
output 	out_data_buffer_62;
output 	out_data_buffer_49;
output 	out_data_buffer_51;
output 	out_data_buffer_50;
output 	out_data_buffer_53;
output 	out_data_buffer_52;
output 	out_data_buffer_55;
output 	out_data_buffer_54;
output 	out_data_buffer_57;
output 	out_data_buffer_56;
output 	out_data_buffer_59;
output 	out_data_buffer_58;
output 	out_data_buffer_61;
output 	out_data_buffer_60;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_buffer_40;
output 	out_data_buffer_41;
output 	out_data_buffer_42;
output 	out_data_buffer_43;
output 	out_data_buffer_44;
output 	out_data_buffer_45;
output 	out_data_buffer_46;
output 	out_data_buffer_47;
output 	out_data_buffer_32;
output 	out_data_buffer_33;
output 	out_data_buffer_34;
output 	out_data_buffer_35;
output 	out_data_buffer_107;
output 	out_data_buffer_86;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_to_out_synchronizer|dreg[0]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_toggle~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \out_data_toggle_flopped~q ;
wire \take_in_data~combout ;
wire \in_data_buffer[68]~q ;
wire \in_data_buffer[48]~q ;
wire \in_data_buffer[62]~q ;
wire \in_data_buffer[49]~q ;
wire \in_data_buffer[51]~q ;
wire \in_data_buffer[50]~q ;
wire \in_data_buffer[53]~q ;
wire \in_data_buffer[52]~q ;
wire \in_data_buffer[55]~q ;
wire \in_data_buffer[54]~q ;
wire \in_data_buffer[57]~q ;
wire \in_data_buffer[56]~q ;
wire \in_data_buffer[59]~q ;
wire \in_data_buffer[58]~q ;
wire \in_data_buffer[61]~q ;
wire \in_data_buffer[60]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \in_data_buffer[40]~q ;
wire \in_data_buffer[41]~q ;
wire \in_data_buffer[42]~q ;
wire \in_data_buffer[43]~q ;
wire \in_data_buffer[44]~q ;
wire \in_data_buffer[45]~q ;
wire \in_data_buffer[46]~q ;
wire \in_data_buffer[47]~q ;
wire \in_data_buffer[32]~q ;
wire \in_data_buffer[33]~q ;
wire \in_data_buffer[34]~q ;
wire \in_data_buffer[35]~q ;
wire \in_data_buffer[107]~q ;
wire \in_data_buffer[86]~q ;


final_project_soc_altera_std_synchronizer_6 out_to_in_synchronizer(
	.reset_n(in_reset),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ),
	.din(\out_data_toggle_flopped~q ),
	.clk(clk_clk));

final_project_soc_altera_std_synchronizer_5 in_to_out_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(out_reset),
	.din(\in_data_toggle~q ),
	.dreg_0(\in_to_out_synchronizer|dreg[0]~q ));

cycloneive_lcell_comb \in_ready~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(in_ready),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h0FF0;
defparam \in_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_data_toggle_flopped~q ),
	.datad(\in_to_out_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[68] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[68]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_68),
	.prn(vcc));
defparam \out_data_buffer[68] .is_wysiwyg = "true";
defparam \out_data_buffer[68] .power_up = "low";

dffeas \out_data_buffer[48] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[48]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_48),
	.prn(vcc));
defparam \out_data_buffer[48] .is_wysiwyg = "true";
defparam \out_data_buffer[48] .power_up = "low";

dffeas \out_data_buffer[62] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[62]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_62),
	.prn(vcc));
defparam \out_data_buffer[62] .is_wysiwyg = "true";
defparam \out_data_buffer[62] .power_up = "low";

dffeas \out_data_buffer[49] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[49]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_49),
	.prn(vcc));
defparam \out_data_buffer[49] .is_wysiwyg = "true";
defparam \out_data_buffer[49] .power_up = "low";

dffeas \out_data_buffer[51] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[51]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_51),
	.prn(vcc));
defparam \out_data_buffer[51] .is_wysiwyg = "true";
defparam \out_data_buffer[51] .power_up = "low";

dffeas \out_data_buffer[50] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[50]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_50),
	.prn(vcc));
defparam \out_data_buffer[50] .is_wysiwyg = "true";
defparam \out_data_buffer[50] .power_up = "low";

dffeas \out_data_buffer[53] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[53]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_53),
	.prn(vcc));
defparam \out_data_buffer[53] .is_wysiwyg = "true";
defparam \out_data_buffer[53] .power_up = "low";

dffeas \out_data_buffer[52] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[52]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_52),
	.prn(vcc));
defparam \out_data_buffer[52] .is_wysiwyg = "true";
defparam \out_data_buffer[52] .power_up = "low";

dffeas \out_data_buffer[55] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[55]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_55),
	.prn(vcc));
defparam \out_data_buffer[55] .is_wysiwyg = "true";
defparam \out_data_buffer[55] .power_up = "low";

dffeas \out_data_buffer[54] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[54]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_54),
	.prn(vcc));
defparam \out_data_buffer[54] .is_wysiwyg = "true";
defparam \out_data_buffer[54] .power_up = "low";

dffeas \out_data_buffer[57] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[57]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_57),
	.prn(vcc));
defparam \out_data_buffer[57] .is_wysiwyg = "true";
defparam \out_data_buffer[57] .power_up = "low";

dffeas \out_data_buffer[56] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[56]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_56),
	.prn(vcc));
defparam \out_data_buffer[56] .is_wysiwyg = "true";
defparam \out_data_buffer[56] .power_up = "low";

dffeas \out_data_buffer[59] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[59]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_59),
	.prn(vcc));
defparam \out_data_buffer[59] .is_wysiwyg = "true";
defparam \out_data_buffer[59] .power_up = "low";

dffeas \out_data_buffer[58] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[58]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_58),
	.prn(vcc));
defparam \out_data_buffer[58] .is_wysiwyg = "true";
defparam \out_data_buffer[58] .power_up = "low";

dffeas \out_data_buffer[61] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[61]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_61),
	.prn(vcc));
defparam \out_data_buffer[61] .is_wysiwyg = "true";
defparam \out_data_buffer[61] .power_up = "low";

dffeas \out_data_buffer[60] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[60]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_60),
	.prn(vcc));
defparam \out_data_buffer[60] .is_wysiwyg = "true";
defparam \out_data_buffer[60] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas \out_data_buffer[40] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[40]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_40),
	.prn(vcc));
defparam \out_data_buffer[40] .is_wysiwyg = "true";
defparam \out_data_buffer[40] .power_up = "low";

dffeas \out_data_buffer[41] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[41]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_41),
	.prn(vcc));
defparam \out_data_buffer[41] .is_wysiwyg = "true";
defparam \out_data_buffer[41] .power_up = "low";

dffeas \out_data_buffer[42] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[42]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_42),
	.prn(vcc));
defparam \out_data_buffer[42] .is_wysiwyg = "true";
defparam \out_data_buffer[42] .power_up = "low";

dffeas \out_data_buffer[43] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[43]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_43),
	.prn(vcc));
defparam \out_data_buffer[43] .is_wysiwyg = "true";
defparam \out_data_buffer[43] .power_up = "low";

dffeas \out_data_buffer[44] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[44]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_44),
	.prn(vcc));
defparam \out_data_buffer[44] .is_wysiwyg = "true";
defparam \out_data_buffer[44] .power_up = "low";

dffeas \out_data_buffer[45] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[45]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_45),
	.prn(vcc));
defparam \out_data_buffer[45] .is_wysiwyg = "true";
defparam \out_data_buffer[45] .power_up = "low";

dffeas \out_data_buffer[46] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[46]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_46),
	.prn(vcc));
defparam \out_data_buffer[46] .is_wysiwyg = "true";
defparam \out_data_buffer[46] .power_up = "low";

dffeas \out_data_buffer[47] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[47]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_47),
	.prn(vcc));
defparam \out_data_buffer[47] .is_wysiwyg = "true";
defparam \out_data_buffer[47] .power_up = "low";

dffeas \out_data_buffer[32] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[32]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_32),
	.prn(vcc));
defparam \out_data_buffer[32] .is_wysiwyg = "true";
defparam \out_data_buffer[32] .power_up = "low";

dffeas \out_data_buffer[33] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[33]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_33),
	.prn(vcc));
defparam \out_data_buffer[33] .is_wysiwyg = "true";
defparam \out_data_buffer[33] .power_up = "low";

dffeas \out_data_buffer[34] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[34]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_34),
	.prn(vcc));
defparam \out_data_buffer[34] .is_wysiwyg = "true";
defparam \out_data_buffer[34] .power_up = "low";

dffeas \out_data_buffer[35] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[35]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_35),
	.prn(vcc));
defparam \out_data_buffer[35] .is_wysiwyg = "true";
defparam \out_data_buffer[35] .power_up = "low";

dffeas \out_data_buffer[107] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[107]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_107),
	.prn(vcc));
defparam \out_data_buffer[107] .is_wysiwyg = "true";
defparam \out_data_buffer[107] .power_up = "low";

dffeas \out_data_buffer[86] (
	.clk(wire_pll7_clk_0),
	.d(\in_data_buffer[86]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_86),
	.prn(vcc));
defparam \out_data_buffer[86] .is_wysiwyg = "true";
defparam \out_data_buffer[86] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(\in_data_toggle~q ),
	.datab(uav_read),
	.datac(src_channel_5),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(\in_to_out_synchronizer|dreg[0]~q ),
	.datab(\out_data_toggle_flopped~q ),
	.datac(last_cycle),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas out_data_toggle_flopped(
	.clk(wire_pll7_clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_toggle_flopped~q ),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb take_in_data(
	.dataa(uav_read),
	.datab(src_channel_5),
	.datac(\in_data_toggle~q ),
	.datad(\out_to_in_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hEFFE;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[68] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[68]~q ),
	.prn(vcc));
defparam \in_data_buffer[68] .is_wysiwyg = "true";
defparam \in_data_buffer[68] .power_up = "low";

dffeas \in_data_buffer[48] (
	.clk(clk_clk),
	.d(in_data[48]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[48]~q ),
	.prn(vcc));
defparam \in_data_buffer[48] .is_wysiwyg = "true";
defparam \in_data_buffer[48] .power_up = "low";

dffeas \in_data_buffer[62] (
	.clk(clk_clk),
	.d(in_data[62]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[62]~q ),
	.prn(vcc));
defparam \in_data_buffer[62] .is_wysiwyg = "true";
defparam \in_data_buffer[62] .power_up = "low";

dffeas \in_data_buffer[49] (
	.clk(clk_clk),
	.d(in_data[49]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[49]~q ),
	.prn(vcc));
defparam \in_data_buffer[49] .is_wysiwyg = "true";
defparam \in_data_buffer[49] .power_up = "low";

dffeas \in_data_buffer[51] (
	.clk(clk_clk),
	.d(in_data[51]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[51]~q ),
	.prn(vcc));
defparam \in_data_buffer[51] .is_wysiwyg = "true";
defparam \in_data_buffer[51] .power_up = "low";

dffeas \in_data_buffer[50] (
	.clk(clk_clk),
	.d(in_data[50]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[50]~q ),
	.prn(vcc));
defparam \in_data_buffer[50] .is_wysiwyg = "true";
defparam \in_data_buffer[50] .power_up = "low";

dffeas \in_data_buffer[53] (
	.clk(clk_clk),
	.d(in_data[53]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[53]~q ),
	.prn(vcc));
defparam \in_data_buffer[53] .is_wysiwyg = "true";
defparam \in_data_buffer[53] .power_up = "low";

dffeas \in_data_buffer[52] (
	.clk(clk_clk),
	.d(in_data[52]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[52]~q ),
	.prn(vcc));
defparam \in_data_buffer[52] .is_wysiwyg = "true";
defparam \in_data_buffer[52] .power_up = "low";

dffeas \in_data_buffer[55] (
	.clk(clk_clk),
	.d(in_data[55]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[55]~q ),
	.prn(vcc));
defparam \in_data_buffer[55] .is_wysiwyg = "true";
defparam \in_data_buffer[55] .power_up = "low";

dffeas \in_data_buffer[54] (
	.clk(clk_clk),
	.d(in_data[54]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[54]~q ),
	.prn(vcc));
defparam \in_data_buffer[54] .is_wysiwyg = "true";
defparam \in_data_buffer[54] .power_up = "low";

dffeas \in_data_buffer[57] (
	.clk(clk_clk),
	.d(in_data[57]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[57]~q ),
	.prn(vcc));
defparam \in_data_buffer[57] .is_wysiwyg = "true";
defparam \in_data_buffer[57] .power_up = "low";

dffeas \in_data_buffer[56] (
	.clk(clk_clk),
	.d(in_data[56]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[56]~q ),
	.prn(vcc));
defparam \in_data_buffer[56] .is_wysiwyg = "true";
defparam \in_data_buffer[56] .power_up = "low";

dffeas \in_data_buffer[59] (
	.clk(clk_clk),
	.d(in_data[59]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[59]~q ),
	.prn(vcc));
defparam \in_data_buffer[59] .is_wysiwyg = "true";
defparam \in_data_buffer[59] .power_up = "low";

dffeas \in_data_buffer[58] (
	.clk(clk_clk),
	.d(in_data[58]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[58]~q ),
	.prn(vcc));
defparam \in_data_buffer[58] .is_wysiwyg = "true";
defparam \in_data_buffer[58] .power_up = "low";

dffeas \in_data_buffer[61] (
	.clk(clk_clk),
	.d(in_data[61]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[61]~q ),
	.prn(vcc));
defparam \in_data_buffer[61] .is_wysiwyg = "true";
defparam \in_data_buffer[61] .power_up = "low";

dffeas \in_data_buffer[60] (
	.clk(clk_clk),
	.d(in_data[60]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[60]~q ),
	.prn(vcc));
defparam \in_data_buffer[60] .is_wysiwyg = "true";
defparam \in_data_buffer[60] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(clk_clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(clk_clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

dffeas \in_data_buffer[40] (
	.clk(clk_clk),
	.d(in_data[40]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[40]~q ),
	.prn(vcc));
defparam \in_data_buffer[40] .is_wysiwyg = "true";
defparam \in_data_buffer[40] .power_up = "low";

dffeas \in_data_buffer[41] (
	.clk(clk_clk),
	.d(in_data[41]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[41]~q ),
	.prn(vcc));
defparam \in_data_buffer[41] .is_wysiwyg = "true";
defparam \in_data_buffer[41] .power_up = "low";

dffeas \in_data_buffer[42] (
	.clk(clk_clk),
	.d(in_data[42]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[42]~q ),
	.prn(vcc));
defparam \in_data_buffer[42] .is_wysiwyg = "true";
defparam \in_data_buffer[42] .power_up = "low";

dffeas \in_data_buffer[43] (
	.clk(clk_clk),
	.d(in_data[43]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[43]~q ),
	.prn(vcc));
defparam \in_data_buffer[43] .is_wysiwyg = "true";
defparam \in_data_buffer[43] .power_up = "low";

dffeas \in_data_buffer[44] (
	.clk(clk_clk),
	.d(in_data[44]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[44]~q ),
	.prn(vcc));
defparam \in_data_buffer[44] .is_wysiwyg = "true";
defparam \in_data_buffer[44] .power_up = "low";

dffeas \in_data_buffer[45] (
	.clk(clk_clk),
	.d(in_data[45]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[45]~q ),
	.prn(vcc));
defparam \in_data_buffer[45] .is_wysiwyg = "true";
defparam \in_data_buffer[45] .power_up = "low";

dffeas \in_data_buffer[46] (
	.clk(clk_clk),
	.d(in_data[46]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[46]~q ),
	.prn(vcc));
defparam \in_data_buffer[46] .is_wysiwyg = "true";
defparam \in_data_buffer[46] .power_up = "low";

dffeas \in_data_buffer[47] (
	.clk(clk_clk),
	.d(in_data[47]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[47]~q ),
	.prn(vcc));
defparam \in_data_buffer[47] .is_wysiwyg = "true";
defparam \in_data_buffer[47] .power_up = "low";

dffeas \in_data_buffer[32] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[32]~q ),
	.prn(vcc));
defparam \in_data_buffer[32] .is_wysiwyg = "true";
defparam \in_data_buffer[32] .power_up = "low";

dffeas \in_data_buffer[33] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[33]~q ),
	.prn(vcc));
defparam \in_data_buffer[33] .is_wysiwyg = "true";
defparam \in_data_buffer[33] .power_up = "low";

dffeas \in_data_buffer[34] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[34]~q ),
	.prn(vcc));
defparam \in_data_buffer[34] .is_wysiwyg = "true";
defparam \in_data_buffer[34] .power_up = "low";

dffeas \in_data_buffer[35] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[35]~q ),
	.prn(vcc));
defparam \in_data_buffer[35] .is_wysiwyg = "true";
defparam \in_data_buffer[35] .power_up = "low";

dffeas \in_data_buffer[107] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[107]~q ),
	.prn(vcc));
defparam \in_data_buffer[107] .is_wysiwyg = "true";
defparam \in_data_buffer[107] .power_up = "low";

dffeas \in_data_buffer[86] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[86]~q ),
	.prn(vcc));
defparam \in_data_buffer[86] .is_wysiwyg = "true";
defparam \in_data_buffer[86] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_5 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_6 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_4 (
	clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_buffer_67,
	in_data_toggle,
	dreg_01,
	take_in_data,
	mem_67_0,
	rp_valid,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_11,
	out_data_13,
	out_data_16,
	out_data_12,
	out_data_5,
	out_data_14,
	out_data_15,
	out_data_21,
	out_data_18,
	out_data_17,
	out_data_31,
	out_data_30,
	out_data_29,
	out_data_28,
	out_data_buffer_31,
	out_data_27,
	out_data_buffer_30,
	out_data_26,
	out_data_buffer_29,
	out_data_25,
	out_data_10,
	out_data_24,
	out_data_9,
	out_data_23,
	out_data_8,
	out_data_22,
	out_data_7,
	out_data_6,
	out_data_20,
	out_data_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
output 	out_data_buffer_67;
output 	in_data_toggle;
output 	dreg_01;
input 	take_in_data;
input 	mem_67_0;
input 	rp_valid;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_11;
input 	out_data_13;
input 	out_data_16;
input 	out_data_12;
input 	out_data_5;
input 	out_data_14;
input 	out_data_15;
input 	out_data_21;
input 	out_data_18;
input 	out_data_17;
input 	out_data_31;
input 	out_data_30;
input 	out_data_29;
input 	out_data_28;
output 	out_data_buffer_31;
input 	out_data_27;
output 	out_data_buffer_30;
input 	out_data_26;
output 	out_data_buffer_29;
input 	out_data_25;
input 	out_data_10;
input 	out_data_24;
input 	out_data_9;
input 	out_data_23;
input 	out_data_8;
input 	out_data_22;
input 	out_data_7;
input 	out_data_6;
input 	out_data_20;
input 	out_data_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_3 clock_xer(
	.clk_0(clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.in_data_toggle1(in_data_toggle),
	.dreg_01(dreg_01),
	.take_in_data(take_in_data),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,mem_67_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_data_31,out_data_30,out_data_29,out_data_28,out_data_27,out_data_26,out_data_25,out_data_24,out_data_23,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,out_data_10,
out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.rp_valid(rp_valid),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_3 (
	clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	out_data_buffer_67,
	in_data_toggle1,
	dreg_01,
	take_in_data,
	in_data,
	rp_valid,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
output 	out_data_buffer_67;
output 	in_data_toggle1;
output 	dreg_01;
input 	take_in_data;
input 	[118:0] in_data;
input 	rp_valid;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \take_in_data~0_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;


final_project_soc_altera_std_synchronizer_8 out_to_in_synchronizer(
	.clk(clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(dreg_01));

final_project_soc_altera_std_synchronizer_7 in_to_out_synchronizer(
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(in_data_toggle1),
	.clk(clk_clk));

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_clk),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas in_data_toggle(
	.clk(clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_clk),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_clk),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(clk_clk),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_clk),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_clk),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_clk),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_clk),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_clk),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_clk),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_clk),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_clk),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_clk),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_clk),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_clk),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_clk),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_clk),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_clk),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_clk),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_clk),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_clk),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_clk),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_clk),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_clk),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(rp_valid),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(take_in_data),
	.cin(gnd),
	.combout(\take_in_data~0_combout ),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hBEFF;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(clk_0),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(take_in_data),
	.datac(rp_valid),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_7 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_8 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_5 (
	clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_valid,
	out_data_buffer_67,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	mem_86_0,
	mem_68_0,
	in_data_toggle,
	dreg_0,
	take_in_data,
	mem_67_0,
	rp_valid,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_21,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_10,
	out_data_buffer_24,
	out_data_buffer_9,
	out_data_buffer_23,
	out_data_buffer_8,
	out_data_buffer_22,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_11,
	out_data_13,
	out_data_16,
	out_data_12,
	out_data_5,
	out_data_14,
	out_data_15,
	out_data_21,
	out_data_18,
	out_data_17,
	out_data_31,
	out_data_30,
	out_data_29,
	out_data_28,
	out_data_27,
	out_data_26,
	out_data_25,
	out_data_10,
	out_data_24,
	out_data_9,
	out_data_23,
	out_data_8,
	out_data_22,
	out_data_7,
	out_data_6,
	out_data_20,
	out_data_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_valid;
output 	out_data_buffer_67;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
input 	mem_86_0;
input 	mem_68_0;
output 	in_data_toggle;
output 	dreg_0;
output 	take_in_data;
input 	mem_67_0;
input 	rp_valid;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_21;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_10;
output 	out_data_buffer_24;
output 	out_data_buffer_9;
output 	out_data_buffer_23;
output 	out_data_buffer_8;
output 	out_data_buffer_22;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_11;
input 	out_data_13;
input 	out_data_16;
input 	out_data_12;
input 	out_data_5;
input 	out_data_14;
input 	out_data_15;
input 	out_data_21;
input 	out_data_18;
input 	out_data_17;
input 	out_data_31;
input 	out_data_30;
input 	out_data_29;
input 	out_data_28;
input 	out_data_27;
input 	out_data_26;
input 	out_data_25;
input 	out_data_10;
input 	out_data_24;
input 	out_data_9;
input 	out_data_23;
input 	out_data_8;
input 	out_data_22;
input 	out_data_7;
input 	out_data_6;
input 	out_data_20;
input 	out_data_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_4 clock_xer(
	.clk_0(clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.in_data_toggle1(in_data_toggle),
	.dreg_0(dreg_0),
	.take_in_data(take_in_data),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,mem_67_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_data_31,out_data_30,out_data_29,out_data_28,out_data_27,out_data_26,out_data_25,out_data_24,out_data_23,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,out_data_10,
out_data_9,out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.rp_valid(rp_valid),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_4 (
	clk_0,
	out_reset,
	in_reset,
	out_valid1,
	out_data_buffer_67,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	mem_86_0,
	mem_68_0,
	in_data_toggle1,
	dreg_0,
	take_in_data,
	in_data,
	rp_valid,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_21,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_10,
	out_data_buffer_24,
	out_data_buffer_9,
	out_data_buffer_23,
	out_data_buffer_8,
	out_data_buffer_22,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_20,
	out_data_buffer_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	out_reset;
input 	in_reset;
output 	out_valid1;
output 	out_data_buffer_67;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
input 	mem_86_0;
input 	mem_68_0;
output 	in_data_toggle1;
output 	dreg_0;
output 	take_in_data;
input 	[118:0] in_data;
input 	rp_valid;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_21;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_10;
output 	out_data_buffer_24;
output 	out_data_buffer_9;
output 	out_data_buffer_23;
output 	out_data_buffer_8;
output 	out_data_buffer_22;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_to_out_synchronizer|dreg[0]~q ;
wire \out_data_toggle_flopped~q ;
wire \take_in_data~1_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;


final_project_soc_altera_std_synchronizer_10 out_to_in_synchronizer(
	.clk(clk_0),
	.reset_n(in_reset),
	.din(\out_data_toggle_flopped~q ),
	.dreg_0(dreg_0));

final_project_soc_altera_std_synchronizer_9 in_to_out_synchronizer(
	.reset_n(out_reset),
	.dreg_0(\in_to_out_synchronizer|dreg[0]~q ),
	.din(in_data_toggle1),
	.clk(clk_clk));

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_data_toggle_flopped~q ),
	.datad(\in_to_out_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_clk),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas in_data_toggle(
	.clk(clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(mem_86_0),
	.datab(mem_68_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(take_in_data),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hEEEE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \out_data_buffer[11] (
	.clk(clk_clk),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_clk),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_clk),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_clk),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_clk),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_clk),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_clk),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_clk),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_clk),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_clk),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_clk),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_clk),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_clk),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_clk),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_clk),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_clk),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_clk),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_clk),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_clk),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_clk),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_clk),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_clk),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_clk),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(\in_to_out_synchronizer|dreg[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_toggle_flopped~q ),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb \take_in_data~1 (
	.dataa(take_in_data),
	.datab(rp_valid),
	.datac(in_data_toggle1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\take_in_data~1_combout ),
	.cout());
defparam \take_in_data~1 .lut_mask = 16'hEFFE;
defparam \take_in_data~1 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(clk_0),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(take_in_data),
	.datac(rp_valid),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[11] (
	.clk(clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_9 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_10 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_6 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_buffer_67,
	mem_used_0,
	mem_107_0,
	out_valid1,
	in_data_toggle,
	dreg_01,
	always0,
	mem_67_0,
	take_in_data,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_11,
	out_payload_13,
	out_payload_16,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_21,
	out_payload_18,
	out_payload_17,
	out_payload_31,
	out_payload_30,
	out_payload_29,
	out_payload_28,
	out_data_buffer_31,
	out_payload_27,
	out_data_buffer_30,
	out_payload_26,
	out_data_buffer_29,
	out_payload_25,
	out_payload_10,
	out_payload_24,
	out_payload_9,
	out_payload_23,
	out_payload_8,
	out_payload_22,
	out_payload_7,
	out_payload_6,
	out_payload_20,
	out_payload_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_toggle_flopped;
output 	dreg_0;
output 	out_valid;
output 	out_data_buffer_67;
input 	mem_used_0;
input 	mem_107_0;
input 	out_valid1;
output 	in_data_toggle;
output 	dreg_01;
input 	always0;
input 	mem_67_0;
output 	take_in_data;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
input 	out_payload_0;
input 	out_payload_1;
input 	out_payload_2;
input 	out_payload_3;
input 	out_payload_4;
input 	out_payload_11;
input 	out_payload_13;
input 	out_payload_16;
input 	out_payload_12;
input 	out_payload_5;
input 	out_payload_14;
input 	out_payload_15;
input 	out_payload_21;
input 	out_payload_18;
input 	out_payload_17;
input 	out_payload_31;
input 	out_payload_30;
input 	out_payload_29;
input 	out_payload_28;
output 	out_data_buffer_31;
input 	out_payload_27;
output 	out_data_buffer_30;
input 	out_payload_26;
output 	out_data_buffer_29;
input 	out_payload_25;
input 	out_payload_10;
input 	out_payload_24;
input 	out_payload_9;
input 	out_payload_23;
input 	out_payload_8;
input 	out_payload_22;
input 	out_payload_7;
input 	out_payload_6;
input 	out_payload_20;
input 	out_payload_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_5 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_data_toggle_flopped1(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.mem_used_0(mem_used_0),
	.mem_107_0(mem_107_0),
	.out_valid2(out_valid1),
	.in_data_toggle1(in_data_toggle),
	.dreg_01(dreg_01),
	.always0(always0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,mem_67_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_payload_31,out_payload_30,out_payload_29,out_payload_28,out_payload_27,out_payload_26,out_payload_25,out_payload_24,out_payload_23,out_payload_22,out_payload_21,out_payload_20,out_payload_19,out_payload_18,out_payload_17,out_payload_16,out_payload_15,
out_payload_14,out_payload_13,out_payload_12,out_payload_11,out_payload_10,out_payload_9,out_payload_8,out_payload_7,out_payload_6,out_payload_5,out_payload_4,out_payload_3,out_payload_2,out_payload_1,out_payload_0}),
	.take_in_data(take_in_data),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_5 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	out_data_buffer_67,
	mem_used_0,
	mem_107_0,
	out_valid2,
	in_data_toggle1,
	dreg_01,
	always0,
	in_data,
	take_in_data,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	out_data_buffer_5,
	out_data_buffer_6,
	out_data_buffer_7,
	out_data_buffer_8,
	out_data_buffer_9,
	out_data_buffer_10,
	out_data_buffer_11,
	out_data_buffer_12,
	out_data_buffer_13,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_16,
	out_data_buffer_17,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
output 	out_data_buffer_67;
input 	mem_used_0;
input 	mem_107_0;
input 	out_valid2;
output 	in_data_toggle1;
output 	dreg_01;
input 	always0;
input 	[118:0] in_data;
output 	take_in_data;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	out_data_buffer_5;
output 	out_data_buffer_6;
output 	out_data_buffer_7;
output 	out_data_buffer_8;
output 	out_data_buffer_9;
output 	out_data_buffer_10;
output 	out_data_buffer_11;
output 	out_data_buffer_12;
output 	out_data_buffer_13;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_16;
output 	out_data_buffer_17;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \take_in_data~1_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;


final_project_soc_altera_std_synchronizer_12 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(out_data_toggle_flopped1),
	.dreg_0(dreg_01));

final_project_soc_altera_std_synchronizer_11 in_to_out_synchronizer(
	.reset_n(out_reset),
	.dreg_0(dreg_0),
	.din(in_data_toggle1),
	.clk(clk_clk));

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(dreg_0),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_clk),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(out_valid2),
	.datab(mem_used_0),
	.datac(mem_107_0),
	.datad(gnd),
	.cin(gnd),
	.combout(take_in_data),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hFEFE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_clk),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_clk),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(clk_clk),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_clk),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_clk),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_clk),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_clk),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_clk),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_clk),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_clk),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_clk),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_clk),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_clk),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_clk),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_clk),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_clk),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_clk),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_clk),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_clk),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_clk),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_clk),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_clk),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_clk),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

cycloneive_lcell_comb \take_in_data~1 (
	.dataa(take_in_data),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(always0),
	.cin(gnd),
	.combout(\take_in_data~1_combout ),
	.cout());
defparam \take_in_data~1 .lut_mask = 16'hBEFF;
defparam \take_in_data~1 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(wire_pll7_clk_0),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(always0),
	.datac(take_in_data),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~1_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_11 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_12 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_handshake_clock_crosser_7 (
	wire_pll7_clk_0,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	out_valid,
	out_data_buffer_67,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	in_data_toggle,
	dreg_0,
	always0,
	mem_67_0,
	take_in_data,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_21,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_10,
	out_data_buffer_24,
	out_data_buffer_9,
	out_data_buffer_23,
	out_data_buffer_8,
	out_data_buffer_22,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_20,
	out_data_buffer_19,
	out_payload_0,
	out_payload_1,
	out_payload_2,
	out_payload_3,
	out_payload_4,
	out_payload_11,
	out_payload_13,
	out_payload_16,
	out_payload_12,
	out_payload_5,
	out_payload_14,
	out_payload_15,
	out_payload_21,
	out_payload_18,
	out_payload_17,
	out_payload_31,
	out_payload_30,
	out_payload_29,
	out_payload_28,
	out_payload_27,
	out_payload_26,
	out_payload_25,
	out_payload_10,
	out_payload_24,
	out_payload_9,
	out_payload_23,
	out_payload_8,
	out_payload_22,
	out_payload_7,
	out_payload_6,
	out_payload_20,
	out_payload_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_valid;
output 	out_data_buffer_67;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	in_data_toggle;
output 	dreg_0;
input 	always0;
input 	mem_67_0;
input 	take_in_data;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_21;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_10;
output 	out_data_buffer_24;
output 	out_data_buffer_9;
output 	out_data_buffer_23;
output 	out_data_buffer_8;
output 	out_data_buffer_22;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
input 	out_payload_0;
input 	out_payload_1;
input 	out_payload_2;
input 	out_payload_3;
input 	out_payload_4;
input 	out_payload_11;
input 	out_payload_13;
input 	out_payload_16;
input 	out_payload_12;
input 	out_payload_5;
input 	out_payload_14;
input 	out_payload_15;
input 	out_payload_21;
input 	out_payload_18;
input 	out_payload_17;
input 	out_payload_31;
input 	out_payload_30;
input 	out_payload_29;
input 	out_payload_28;
input 	out_payload_27;
input 	out_payload_26;
input 	out_payload_25;
input 	out_payload_10;
input 	out_payload_24;
input 	out_payload_9;
input 	out_payload_23;
input 	out_payload_8;
input 	out_payload_22;
input 	out_payload_7;
input 	out_payload_6;
input 	out_payload_20;
input 	out_payload_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_avalon_st_clock_crosser_6 clock_xer(
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.out_reset(r_sync_rst),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.out_valid1(out_valid),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_1(out_data_buffer_1),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_4(out_data_buffer_4),
	.in_data_toggle1(in_data_toggle),
	.dreg_0(dreg_0),
	.always0(always0),
	.in_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,mem_67_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,out_payload_31,out_payload_30,out_payload_29,out_payload_28,out_payload_27,out_payload_26,out_payload_25,out_payload_24,out_payload_23,out_payload_22,out_payload_21,out_payload_20,out_payload_19,out_payload_18,out_payload_17,out_payload_16,out_payload_15,
out_payload_14,out_payload_13,out_payload_12,out_payload_11,out_payload_10,out_payload_9,out_payload_8,out_payload_7,out_payload_6,out_payload_5,out_payload_4,out_payload_3,out_payload_2,out_payload_1,out_payload_0}),
	.take_in_data(take_in_data),
	.out_data_buffer_11(out_data_buffer_11),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_14(out_data_buffer_14),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_21(out_data_buffer_21),
	.out_data_buffer_18(out_data_buffer_18),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_31(out_data_buffer_31),
	.out_data_buffer_30(out_data_buffer_30),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_28(out_data_buffer_28),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_26(out_data_buffer_26),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_10(out_data_buffer_10),
	.out_data_buffer_24(out_data_buffer_24),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_8(out_data_buffer_8),
	.out_data_buffer_22(out_data_buffer_22),
	.out_data_buffer_7(out_data_buffer_7),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_19(out_data_buffer_19),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_6 (
	wire_pll7_clk_0,
	out_reset,
	in_reset,
	out_valid1,
	out_data_buffer_67,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_3,
	out_data_buffer_4,
	in_data_toggle1,
	dreg_0,
	always0,
	in_data,
	take_in_data,
	out_data_buffer_11,
	out_data_buffer_13,
	out_data_buffer_16,
	out_data_buffer_12,
	out_data_buffer_5,
	out_data_buffer_14,
	out_data_buffer_15,
	out_data_buffer_21,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_31,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_10,
	out_data_buffer_24,
	out_data_buffer_9,
	out_data_buffer_23,
	out_data_buffer_8,
	out_data_buffer_22,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_20,
	out_data_buffer_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	out_reset;
input 	in_reset;
output 	out_valid1;
output 	out_data_buffer_67;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_3;
output 	out_data_buffer_4;
output 	in_data_toggle1;
output 	dreg_0;
input 	always0;
input 	[118:0] in_data;
input 	take_in_data;
output 	out_data_buffer_11;
output 	out_data_buffer_13;
output 	out_data_buffer_16;
output 	out_data_buffer_12;
output 	out_data_buffer_5;
output 	out_data_buffer_14;
output 	out_data_buffer_15;
output 	out_data_buffer_21;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_31;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_10;
output 	out_data_buffer_24;
output 	out_data_buffer_9;
output 	out_data_buffer_23;
output 	out_data_buffer_8;
output 	out_data_buffer_22;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_to_out_synchronizer|dreg[0]~q ;
wire \out_data_toggle_flopped~q ;
wire \take_in_data~0_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;


final_project_soc_altera_std_synchronizer_14 out_to_in_synchronizer(
	.clk(wire_pll7_clk_0),
	.reset_n(in_reset),
	.din(\out_data_toggle_flopped~q ),
	.dreg_0(dreg_0));

final_project_soc_altera_std_synchronizer_13 in_to_out_synchronizer(
	.reset_n(out_reset),
	.dreg_0(\in_to_out_synchronizer|dreg[0]~q ),
	.din(in_data_toggle1),
	.clk(clk_clk));

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_data_toggle_flopped~q ),
	.datad(\in_to_out_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_clk),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_clk),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_clk),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_clk),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(clk_clk),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_clk),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas in_data_toggle(
	.clk(wire_pll7_clk_0),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(clk_clk),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_clk),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_clk),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_clk),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_clk),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_clk),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_clk),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_clk),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_clk),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_clk),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_clk),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_clk),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_clk),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_clk),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_clk),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_clk),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_clk),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_clk),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_clk),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_clk),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_clk),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_clk),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_clk),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_clk),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_clk),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_clk),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_clk),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(clk_clk),
	.d(\in_to_out_synchronizer|dreg[0]~q ),
	.asdata(vcc),
	.clrn(!out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_toggle_flopped~q ),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(always0),
	.datab(take_in_data),
	.datac(in_data_toggle1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\take_in_data~0_combout ),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hEFFE;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(wire_pll7_clk_0),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(wire_pll7_clk_0),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(wire_pll7_clk_0),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(wire_pll7_clk_0),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(wire_pll7_clk_0),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(wire_pll7_clk_0),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(always0),
	.datac(take_in_data),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hBEFF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[11] (
	.clk(wire_pll7_clk_0),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(wire_pll7_clk_0),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(wire_pll7_clk_0),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(wire_pll7_clk_0),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(wire_pll7_clk_0),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(wire_pll7_clk_0),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(wire_pll7_clk_0),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(wire_pll7_clk_0),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(wire_pll7_clk_0),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(wire_pll7_clk_0),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(wire_pll7_clk_0),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(wire_pll7_clk_0),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(wire_pll7_clk_0),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(wire_pll7_clk_0),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(wire_pll7_clk_0),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(wire_pll7_clk_0),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(wire_pll7_clk_0),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(wire_pll7_clk_0),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(wire_pll7_clk_0),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(wire_pll7_clk_0),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(wire_pll7_clk_0),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(wire_pll7_clk_0),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(wire_pll7_clk_0),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(wire_pll7_clk_0),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(wire_pll7_clk_0),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(wire_pll7_clk_0),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(wire_pll7_clk_0),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~0_combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_13 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_14 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_avalon_st_clock_crosser_7 (
	W_alu_result_4,
	in_data,
	clk_0,
	cp_valid,
	in_reset,
	out_reset,
	Equal3,
	take_in_data1,
	saved_grant_0,
	out_data_buffer_3,
	out_data_buffer_38,
	out_data_buffer_39,
	out_data_toggle_flopped1,
	dreg_0,
	out_valid1,
	out_data_buffer_67,
	out_data_buffer_31,
	out_data_buffer_107,
	mem_used_0,
	out_data_buffer_66,
	out_data_buffer_68,
	out_data_buffer_30,
	out_data_buffer_29,
	out_data_buffer_28,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_27,
	out_data_buffer_26,
	out_data_buffer_25,
	out_data_buffer_24,
	out_data_buffer_23,
	out_data_buffer_22,
	out_data_buffer_21,
	out_data_buffer_20,
	out_data_buffer_19,
	out_data_buffer_18,
	out_data_buffer_17,
	out_data_buffer_16,
	out_data_buffer_15,
	out_data_buffer_14,
	out_data_buffer_13,
	out_data_buffer_12,
	out_data_buffer_11,
	out_data_buffer_10,
	out_data_buffer_9,
	out_data_buffer_8,
	out_data_buffer_7,
	out_data_buffer_6,
	out_data_buffer_5,
	out_data_buffer_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	[118:0] in_data;
input 	clk_0;
input 	cp_valid;
input 	in_reset;
input 	out_reset;
input 	Equal3;
output 	take_in_data1;
input 	saved_grant_0;
output 	out_data_buffer_3;
output 	out_data_buffer_38;
output 	out_data_buffer_39;
output 	out_data_toggle_flopped1;
output 	dreg_0;
output 	out_valid1;
output 	out_data_buffer_67;
output 	out_data_buffer_31;
output 	out_data_buffer_107;
input 	mem_used_0;
output 	out_data_buffer_66;
output 	out_data_buffer_68;
output 	out_data_buffer_30;
output 	out_data_buffer_29;
output 	out_data_buffer_28;
output 	out_data_buffer_0;
output 	out_data_buffer_1;
output 	out_data_buffer_2;
output 	out_data_buffer_27;
output 	out_data_buffer_26;
output 	out_data_buffer_25;
output 	out_data_buffer_24;
output 	out_data_buffer_23;
output 	out_data_buffer_22;
output 	out_data_buffer_21;
output 	out_data_buffer_20;
output 	out_data_buffer_19;
output 	out_data_buffer_18;
output 	out_data_buffer_17;
output 	out_data_buffer_16;
output 	out_data_buffer_15;
output 	out_data_buffer_14;
output 	out_data_buffer_13;
output 	out_data_buffer_12;
output 	out_data_buffer_11;
output 	out_data_buffer_10;
output 	out_data_buffer_9;
output 	out_data_buffer_8;
output 	out_data_buffer_7;
output 	out_data_buffer_6;
output 	out_data_buffer_5;
output 	out_data_buffer_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_to_in_synchronizer|dreg[0]~q ;
wire \in_data_toggle~0_combout ;
wire \in_data_toggle~q ;
wire \take_in_data~combout ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[38]~q ;
wire \in_data_buffer[39]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \in_data_buffer[67]~q ;
wire \in_data_buffer[31]~q ;
wire \in_data_buffer[107]~q ;
wire \in_data_buffer[66]~q ;
wire \in_data_buffer[68]~q ;
wire \in_data_buffer[30]~q ;
wire \in_data_buffer[29]~q ;
wire \in_data_buffer[28]~q ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[27]~q ;
wire \in_data_buffer[26]~q ;
wire \in_data_buffer[25]~q ;
wire \in_data_buffer[24]~q ;
wire \in_data_buffer[23]~q ;
wire \in_data_buffer[22]~q ;
wire \in_data_buffer[21]~q ;
wire \in_data_buffer[20]~q ;
wire \in_data_buffer[19]~q ;
wire \in_data_buffer[18]~q ;
wire \in_data_buffer[17]~q ;
wire \in_data_buffer[16]~q ;
wire \in_data_buffer[15]~q ;
wire \in_data_buffer[14]~q ;
wire \in_data_buffer[13]~q ;
wire \in_data_buffer[12]~q ;
wire \in_data_buffer[11]~q ;
wire \in_data_buffer[10]~q ;
wire \in_data_buffer[9]~q ;
wire \in_data_buffer[8]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[4]~q ;


final_project_soc_altera_std_synchronizer_16 out_to_in_synchronizer(
	.reset_n(in_reset),
	.dreg_0(\out_to_in_synchronizer|dreg[0]~q ),
	.din(out_data_toggle_flopped1),
	.clk(clk_clk));

final_project_soc_altera_std_synchronizer_15 in_to_out_synchronizer(
	.clk(clk_0),
	.reset_n(out_reset),
	.din(\in_data_toggle~q ),
	.dreg_0(dreg_0));

cycloneive_lcell_comb \take_in_data~0 (
	.dataa(Equal3),
	.datab(\in_data_toggle~q ),
	.datac(\out_to_in_synchronizer|dreg[0]~q ),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(take_in_data1),
	.cout());
defparam \take_in_data~0 .lut_mask = 16'hBEFF;
defparam \take_in_data~0 .sum_lutc_input = "datac";

dffeas \out_data_buffer[3] (
	.clk(clk_0),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_3),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[38] (
	.clk(clk_0),
	.d(\in_data_buffer[38]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_38),
	.prn(vcc));
defparam \out_data_buffer[38] .is_wysiwyg = "true";
defparam \out_data_buffer[38] .power_up = "low";

dffeas \out_data_buffer[39] (
	.clk(clk_0),
	.d(\in_data_buffer[39]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_39),
	.prn(vcc));
defparam \out_data_buffer[39] .is_wysiwyg = "true";
defparam \out_data_buffer[39] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(clk_0),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_toggle_flopped1),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

cycloneive_lcell_comb out_valid(
	.dataa(gnd),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_0),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'h0FF0;
defparam out_valid.sum_lutc_input = "datac";

dffeas \out_data_buffer[67] (
	.clk(clk_0),
	.d(\in_data_buffer[67]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_67),
	.prn(vcc));
defparam \out_data_buffer[67] .is_wysiwyg = "true";
defparam \out_data_buffer[67] .power_up = "low";

dffeas \out_data_buffer[31] (
	.clk(clk_0),
	.d(\in_data_buffer[31]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_31),
	.prn(vcc));
defparam \out_data_buffer[31] .is_wysiwyg = "true";
defparam \out_data_buffer[31] .power_up = "low";

dffeas \out_data_buffer[107] (
	.clk(clk_0),
	.d(\in_data_buffer[107]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_107),
	.prn(vcc));
defparam \out_data_buffer[107] .is_wysiwyg = "true";
defparam \out_data_buffer[107] .power_up = "low";

dffeas \out_data_buffer[66] (
	.clk(clk_0),
	.d(\in_data_buffer[66]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_66),
	.prn(vcc));
defparam \out_data_buffer[66] .is_wysiwyg = "true";
defparam \out_data_buffer[66] .power_up = "low";

dffeas \out_data_buffer[68] (
	.clk(clk_0),
	.d(\in_data_buffer[68]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_68),
	.prn(vcc));
defparam \out_data_buffer[68] .is_wysiwyg = "true";
defparam \out_data_buffer[68] .power_up = "low";

dffeas \out_data_buffer[30] (
	.clk(clk_0),
	.d(\in_data_buffer[30]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_30),
	.prn(vcc));
defparam \out_data_buffer[30] .is_wysiwyg = "true";
defparam \out_data_buffer[30] .power_up = "low";

dffeas \out_data_buffer[29] (
	.clk(clk_0),
	.d(\in_data_buffer[29]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_29),
	.prn(vcc));
defparam \out_data_buffer[29] .is_wysiwyg = "true";
defparam \out_data_buffer[29] .power_up = "low";

dffeas \out_data_buffer[28] (
	.clk(clk_0),
	.d(\in_data_buffer[28]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_28),
	.prn(vcc));
defparam \out_data_buffer[28] .is_wysiwyg = "true";
defparam \out_data_buffer[28] .power_up = "low";

dffeas \out_data_buffer[0] (
	.clk(clk_0),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_0),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(clk_0),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_1),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(clk_0),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_2),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[27] (
	.clk(clk_0),
	.d(\in_data_buffer[27]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_27),
	.prn(vcc));
defparam \out_data_buffer[27] .is_wysiwyg = "true";
defparam \out_data_buffer[27] .power_up = "low";

dffeas \out_data_buffer[26] (
	.clk(clk_0),
	.d(\in_data_buffer[26]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_26),
	.prn(vcc));
defparam \out_data_buffer[26] .is_wysiwyg = "true";
defparam \out_data_buffer[26] .power_up = "low";

dffeas \out_data_buffer[25] (
	.clk(clk_0),
	.d(\in_data_buffer[25]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_25),
	.prn(vcc));
defparam \out_data_buffer[25] .is_wysiwyg = "true";
defparam \out_data_buffer[25] .power_up = "low";

dffeas \out_data_buffer[24] (
	.clk(clk_0),
	.d(\in_data_buffer[24]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_24),
	.prn(vcc));
defparam \out_data_buffer[24] .is_wysiwyg = "true";
defparam \out_data_buffer[24] .power_up = "low";

dffeas \out_data_buffer[23] (
	.clk(clk_0),
	.d(\in_data_buffer[23]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_23),
	.prn(vcc));
defparam \out_data_buffer[23] .is_wysiwyg = "true";
defparam \out_data_buffer[23] .power_up = "low";

dffeas \out_data_buffer[22] (
	.clk(clk_0),
	.d(\in_data_buffer[22]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_22),
	.prn(vcc));
defparam \out_data_buffer[22] .is_wysiwyg = "true";
defparam \out_data_buffer[22] .power_up = "low";

dffeas \out_data_buffer[21] (
	.clk(clk_0),
	.d(\in_data_buffer[21]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_21),
	.prn(vcc));
defparam \out_data_buffer[21] .is_wysiwyg = "true";
defparam \out_data_buffer[21] .power_up = "low";

dffeas \out_data_buffer[20] (
	.clk(clk_0),
	.d(\in_data_buffer[20]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_20),
	.prn(vcc));
defparam \out_data_buffer[20] .is_wysiwyg = "true";
defparam \out_data_buffer[20] .power_up = "low";

dffeas \out_data_buffer[19] (
	.clk(clk_0),
	.d(\in_data_buffer[19]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_19),
	.prn(vcc));
defparam \out_data_buffer[19] .is_wysiwyg = "true";
defparam \out_data_buffer[19] .power_up = "low";

dffeas \out_data_buffer[18] (
	.clk(clk_0),
	.d(\in_data_buffer[18]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_18),
	.prn(vcc));
defparam \out_data_buffer[18] .is_wysiwyg = "true";
defparam \out_data_buffer[18] .power_up = "low";

dffeas \out_data_buffer[17] (
	.clk(clk_0),
	.d(\in_data_buffer[17]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_17),
	.prn(vcc));
defparam \out_data_buffer[17] .is_wysiwyg = "true";
defparam \out_data_buffer[17] .power_up = "low";

dffeas \out_data_buffer[16] (
	.clk(clk_0),
	.d(\in_data_buffer[16]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_16),
	.prn(vcc));
defparam \out_data_buffer[16] .is_wysiwyg = "true";
defparam \out_data_buffer[16] .power_up = "low";

dffeas \out_data_buffer[15] (
	.clk(clk_0),
	.d(\in_data_buffer[15]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_15),
	.prn(vcc));
defparam \out_data_buffer[15] .is_wysiwyg = "true";
defparam \out_data_buffer[15] .power_up = "low";

dffeas \out_data_buffer[14] (
	.clk(clk_0),
	.d(\in_data_buffer[14]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_14),
	.prn(vcc));
defparam \out_data_buffer[14] .is_wysiwyg = "true";
defparam \out_data_buffer[14] .power_up = "low";

dffeas \out_data_buffer[13] (
	.clk(clk_0),
	.d(\in_data_buffer[13]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_13),
	.prn(vcc));
defparam \out_data_buffer[13] .is_wysiwyg = "true";
defparam \out_data_buffer[13] .power_up = "low";

dffeas \out_data_buffer[12] (
	.clk(clk_0),
	.d(\in_data_buffer[12]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_12),
	.prn(vcc));
defparam \out_data_buffer[12] .is_wysiwyg = "true";
defparam \out_data_buffer[12] .power_up = "low";

dffeas \out_data_buffer[11] (
	.clk(clk_0),
	.d(\in_data_buffer[11]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_11),
	.prn(vcc));
defparam \out_data_buffer[11] .is_wysiwyg = "true";
defparam \out_data_buffer[11] .power_up = "low";

dffeas \out_data_buffer[10] (
	.clk(clk_0),
	.d(\in_data_buffer[10]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_10),
	.prn(vcc));
defparam \out_data_buffer[10] .is_wysiwyg = "true";
defparam \out_data_buffer[10] .power_up = "low";

dffeas \out_data_buffer[9] (
	.clk(clk_0),
	.d(\in_data_buffer[9]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_9),
	.prn(vcc));
defparam \out_data_buffer[9] .is_wysiwyg = "true";
defparam \out_data_buffer[9] .power_up = "low";

dffeas \out_data_buffer[8] (
	.clk(clk_0),
	.d(\in_data_buffer[8]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_8),
	.prn(vcc));
defparam \out_data_buffer[8] .is_wysiwyg = "true";
defparam \out_data_buffer[8] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(clk_0),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_7),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(clk_0),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_6),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(clk_0),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_5),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(clk_0),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(out_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_buffer_4),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

cycloneive_lcell_comb \in_data_toggle~0 (
	.dataa(gnd),
	.datab(\in_data_toggle~q ),
	.datac(cp_valid),
	.datad(take_in_data1),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hC33C;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_data_toggle~q ),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

cycloneive_lcell_comb take_in_data(
	.dataa(cp_valid),
	.datab(take_in_data1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hEEEE;
defparam take_in_data.sum_lutc_input = "datac";

dffeas \in_data_buffer[3] (
	.clk(clk_clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[38] (
	.clk(clk_clk),
	.d(in_data[38]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[38]~q ),
	.prn(vcc));
defparam \in_data_buffer[38] .is_wysiwyg = "true";
defparam \in_data_buffer[38] .power_up = "low";

dffeas \in_data_buffer[39] (
	.clk(clk_clk),
	.d(in_data[39]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[39]~q ),
	.prn(vcc));
defparam \in_data_buffer[39] .is_wysiwyg = "true";
defparam \in_data_buffer[39] .power_up = "low";

cycloneive_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(dreg_0),
	.datab(out_data_toggle_flopped1),
	.datac(saved_grant_0),
	.datad(mem_used_0),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hEFFE;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

dffeas \in_data_buffer[67] (
	.clk(clk_clk),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[67]~q ),
	.prn(vcc));
defparam \in_data_buffer[67] .is_wysiwyg = "true";
defparam \in_data_buffer[67] .power_up = "low";

dffeas \in_data_buffer[31] (
	.clk(clk_clk),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[31]~q ),
	.prn(vcc));
defparam \in_data_buffer[31] .is_wysiwyg = "true";
defparam \in_data_buffer[31] .power_up = "low";

dffeas \in_data_buffer[107] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[107]~q ),
	.prn(vcc));
defparam \in_data_buffer[107] .is_wysiwyg = "true";
defparam \in_data_buffer[107] .power_up = "low";

dffeas \in_data_buffer[66] (
	.clk(clk_clk),
	.d(in_data[67]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[66]~q ),
	.prn(vcc));
defparam \in_data_buffer[66] .is_wysiwyg = "true";
defparam \in_data_buffer[66] .power_up = "low";

dffeas \in_data_buffer[68] (
	.clk(clk_clk),
	.d(in_data[68]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[68]~q ),
	.prn(vcc));
defparam \in_data_buffer[68] .is_wysiwyg = "true";
defparam \in_data_buffer[68] .power_up = "low";

dffeas \in_data_buffer[30] (
	.clk(clk_clk),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[30]~q ),
	.prn(vcc));
defparam \in_data_buffer[30] .is_wysiwyg = "true";
defparam \in_data_buffer[30] .power_up = "low";

dffeas \in_data_buffer[29] (
	.clk(clk_clk),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[29]~q ),
	.prn(vcc));
defparam \in_data_buffer[29] .is_wysiwyg = "true";
defparam \in_data_buffer[29] .power_up = "low";

dffeas \in_data_buffer[28] (
	.clk(clk_clk),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[28]~q ),
	.prn(vcc));
defparam \in_data_buffer[28] .is_wysiwyg = "true";
defparam \in_data_buffer[28] .power_up = "low";

dffeas \in_data_buffer[0] (
	.clk(clk_clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[27] (
	.clk(clk_clk),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[27]~q ),
	.prn(vcc));
defparam \in_data_buffer[27] .is_wysiwyg = "true";
defparam \in_data_buffer[27] .power_up = "low";

dffeas \in_data_buffer[26] (
	.clk(clk_clk),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[26]~q ),
	.prn(vcc));
defparam \in_data_buffer[26] .is_wysiwyg = "true";
defparam \in_data_buffer[26] .power_up = "low";

dffeas \in_data_buffer[25] (
	.clk(clk_clk),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[25]~q ),
	.prn(vcc));
defparam \in_data_buffer[25] .is_wysiwyg = "true";
defparam \in_data_buffer[25] .power_up = "low";

dffeas \in_data_buffer[24] (
	.clk(clk_clk),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[24]~q ),
	.prn(vcc));
defparam \in_data_buffer[24] .is_wysiwyg = "true";
defparam \in_data_buffer[24] .power_up = "low";

dffeas \in_data_buffer[23] (
	.clk(clk_clk),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[23]~q ),
	.prn(vcc));
defparam \in_data_buffer[23] .is_wysiwyg = "true";
defparam \in_data_buffer[23] .power_up = "low";

dffeas \in_data_buffer[22] (
	.clk(clk_clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[22]~q ),
	.prn(vcc));
defparam \in_data_buffer[22] .is_wysiwyg = "true";
defparam \in_data_buffer[22] .power_up = "low";

dffeas \in_data_buffer[21] (
	.clk(clk_clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[21]~q ),
	.prn(vcc));
defparam \in_data_buffer[21] .is_wysiwyg = "true";
defparam \in_data_buffer[21] .power_up = "low";

dffeas \in_data_buffer[20] (
	.clk(clk_clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[20]~q ),
	.prn(vcc));
defparam \in_data_buffer[20] .is_wysiwyg = "true";
defparam \in_data_buffer[20] .power_up = "low";

dffeas \in_data_buffer[19] (
	.clk(clk_clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[19]~q ),
	.prn(vcc));
defparam \in_data_buffer[19] .is_wysiwyg = "true";
defparam \in_data_buffer[19] .power_up = "low";

dffeas \in_data_buffer[18] (
	.clk(clk_clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[18]~q ),
	.prn(vcc));
defparam \in_data_buffer[18] .is_wysiwyg = "true";
defparam \in_data_buffer[18] .power_up = "low";

dffeas \in_data_buffer[17] (
	.clk(clk_clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[17]~q ),
	.prn(vcc));
defparam \in_data_buffer[17] .is_wysiwyg = "true";
defparam \in_data_buffer[17] .power_up = "low";

dffeas \in_data_buffer[16] (
	.clk(clk_clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[16]~q ),
	.prn(vcc));
defparam \in_data_buffer[16] .is_wysiwyg = "true";
defparam \in_data_buffer[16] .power_up = "low";

dffeas \in_data_buffer[15] (
	.clk(clk_clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[15]~q ),
	.prn(vcc));
defparam \in_data_buffer[15] .is_wysiwyg = "true";
defparam \in_data_buffer[15] .power_up = "low";

dffeas \in_data_buffer[14] (
	.clk(clk_clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[14]~q ),
	.prn(vcc));
defparam \in_data_buffer[14] .is_wysiwyg = "true";
defparam \in_data_buffer[14] .power_up = "low";

dffeas \in_data_buffer[13] (
	.clk(clk_clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[13]~q ),
	.prn(vcc));
defparam \in_data_buffer[13] .is_wysiwyg = "true";
defparam \in_data_buffer[13] .power_up = "low";

dffeas \in_data_buffer[12] (
	.clk(clk_clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[12]~q ),
	.prn(vcc));
defparam \in_data_buffer[12] .is_wysiwyg = "true";
defparam \in_data_buffer[12] .power_up = "low";

dffeas \in_data_buffer[11] (
	.clk(clk_clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[11]~q ),
	.prn(vcc));
defparam \in_data_buffer[11] .is_wysiwyg = "true";
defparam \in_data_buffer[11] .power_up = "low";

dffeas \in_data_buffer[10] (
	.clk(clk_clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[10]~q ),
	.prn(vcc));
defparam \in_data_buffer[10] .is_wysiwyg = "true";
defparam \in_data_buffer[10] .power_up = "low";

dffeas \in_data_buffer[9] (
	.clk(clk_clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[9]~q ),
	.prn(vcc));
defparam \in_data_buffer[9] .is_wysiwyg = "true";
defparam \in_data_buffer[9] .power_up = "low";

dffeas \in_data_buffer[8] (
	.clk(clk_clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[8]~q ),
	.prn(vcc));
defparam \in_data_buffer[8] .is_wysiwyg = "true";
defparam \in_data_buffer[8] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_15 (
	clk,
	reset_n,
	din,
	dreg_0)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	din;
output 	dreg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_16 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_merlin_master_agent (
	d_read,
	d_write,
	read_accepted,
	write_accepted,
	cp_valid1)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	d_write;
input 	read_accepted;
input 	write_accepted;
output 	cp_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb cp_valid(
	.dataa(d_read),
	.datab(d_write),
	.datac(read_accepted),
	.datad(write_accepted),
	.cin(gnd),
	.combout(cp_valid1),
	.cout());
defparam cp_valid.lut_mask = 16'hEFFF;
defparam cp_valid.sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_master_agent_1 (
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	mem_67_04,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src_payload,
	src_payload1,
	out_valid,
	out_valid1,
	WideOr1,
	out_data_buffer_67,
	out_data_buffer_671,
	av_readdatavalid)/* synthesis synthesis_greybox=1 */;
input 	mem_67_0;
input 	mem_67_01;
input 	mem_67_02;
input 	mem_67_03;
input 	mem_67_04;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	src_payload;
input 	src_payload1;
input 	out_valid;
input 	out_valid1;
input 	WideOr1;
input 	out_data_buffer_67;
input 	out_data_buffer_671;
output 	av_readdatavalid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdatavalid~0_combout ;
wire \av_readdatavalid~1_combout ;
wire \av_readdatavalid~2_combout ;
wire \av_readdatavalid~3_combout ;


cycloneive_lcell_comb \av_readdatavalid~4 (
	.dataa(WideOr1),
	.datab(\av_readdatavalid~0_combout ),
	.datac(\av_readdatavalid~1_combout ),
	.datad(\av_readdatavalid~3_combout ),
	.cin(gnd),
	.combout(av_readdatavalid),
	.cout());
defparam \av_readdatavalid~4 .lut_mask = 16'hFFFE;
defparam \av_readdatavalid~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdatavalid~0 (
	.dataa(src1_valid),
	.datab(mem_67_0),
	.datac(src1_valid1),
	.datad(mem_67_02),
	.cin(gnd),
	.combout(\av_readdatavalid~0_combout ),
	.cout());
defparam \av_readdatavalid~0 .lut_mask = 16'h7FFF;
defparam \av_readdatavalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdatavalid~1 (
	.dataa(src1_valid2),
	.datab(mem_67_04),
	.datac(src_payload1),
	.datad(mem_67_01),
	.cin(gnd),
	.combout(\av_readdatavalid~1_combout ),
	.cout());
defparam \av_readdatavalid~1 .lut_mask = 16'h7FFF;
defparam \av_readdatavalid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdatavalid~2 (
	.dataa(out_valid),
	.datab(out_data_buffer_67),
	.datac(out_valid1),
	.datad(out_data_buffer_671),
	.cin(gnd),
	.combout(\av_readdatavalid~2_combout ),
	.cout());
defparam \av_readdatavalid~2 .lut_mask = 16'h7FFF;
defparam \av_readdatavalid~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdatavalid~3 (
	.dataa(\av_readdatavalid~2_combout ),
	.datab(gnd),
	.datac(src_payload),
	.datad(mem_67_03),
	.cin(gnd),
	.combout(\av_readdatavalid~3_combout ),
	.cout());
defparam \av_readdatavalid~3 .lut_mask = 16'hAFFF;
defparam \av_readdatavalid~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_master_translator (
	d_read,
	d_write,
	read_accepted1,
	write_accepted1,
	cp_valid,
	uav_write,
	reset,
	uav_read,
	rst1,
	WideOr0,
	WideOr01,
	av_waitrequest,
	av_ld_getting_data,
	clk)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	d_write;
output 	read_accepted1;
output 	write_accepted1;
input 	cp_valid;
output 	uav_write;
input 	reset;
output 	uav_read;
input 	rst1;
input 	WideOr0;
input 	WideOr01;
output 	av_waitrequest;
input 	av_ld_getting_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write_accepted~0_combout ;
wire \read_accepted~0_combout ;
wire \write_accepted~1_combout ;
wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;
wire \av_waitrequest~0_combout ;
wire \av_waitrequest~1_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

cycloneive_lcell_comb \uav_write~0 (
	.dataa(d_write),
	.datab(gnd),
	.datac(gnd),
	.datad(write_accepted1),
	.cin(gnd),
	.combout(uav_write),
	.cout());
defparam \uav_write~0 .lut_mask = 16'hAAFF;
defparam \uav_write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \uav_read~0 (
	.dataa(d_read),
	.datab(gnd),
	.datac(gnd),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read),
	.cout());
defparam \uav_read~0 .lut_mask = 16'hAAFF;
defparam \uav_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~2 (
	.dataa(d_read),
	.datab(d_write),
	.datac(av_ld_getting_data),
	.datad(\av_waitrequest~1_combout ),
	.cin(gnd),
	.combout(av_waitrequest),
	.cout());
defparam \av_waitrequest~2 .lut_mask = 16'h27FF;
defparam \av_waitrequest~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_accepted~0 (
	.dataa(rst1),
	.datab(WideOr0),
	.datac(WideOr01),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_accepted~0_combout ),
	.cout());
defparam \write_accepted~0 .lut_mask = 16'hFEFE;
defparam \write_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(read_accepted1),
	.datab(d_read),
	.datac(\write_accepted~0_combout ),
	.datad(av_ld_getting_data),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hFEFF;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_accepted~1 (
	.dataa(av_waitrequest),
	.datab(write_accepted1),
	.datac(d_write),
	.datad(\write_accepted~0_combout ),
	.cin(gnd),
	.combout(\write_accepted~1_combout ),
	.cout());
defparam \write_accepted~1 .lut_mask = 16'hFFFE;
defparam \write_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \end_begintransfer~0 (
	.dataa(cp_valid),
	.datab(\end_begintransfer~q ),
	.datac(gnd),
	.datad(\write_accepted~0_combout ),
	.cin(gnd),
	.combout(\end_begintransfer~0_combout ),
	.cout());
defparam \end_begintransfer~0 .lut_mask = 16'hEEFF;
defparam \end_begintransfer~0 .sum_lutc_input = "datac";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(\end_begintransfer~q ),
	.datab(WideOr0),
	.datac(WideOr01),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFEFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~1 (
	.dataa(rst1),
	.datab(write_accepted1),
	.datac(\av_waitrequest~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest~1_combout ),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'hFEFE;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_master_translator_1 (
	saved_grant_1,
	F_pc_5,
	i_read,
	read_accepted1,
	uav_read1,
	F_pc_2,
	mem_used_1,
	reset,
	rst1,
	waitrequest,
	mem_used_11,
	mem_used_12,
	waitrequest1,
	mem_used_13,
	Equal1,
	wait_latency_counter_1,
	av_readdatavalid,
	src_valid,
	Equal0,
	src_channel_6,
	mem,
	Equal6,
	Equal2,
	take_in_data,
	saved_grant_11,
	Equal5,
	saved_grant_12,
	src_channel_5,
	in_ready,
	clk)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_1;
input 	F_pc_5;
input 	i_read;
output 	read_accepted1;
output 	uav_read1;
input 	F_pc_2;
input 	mem_used_1;
input 	reset;
input 	rst1;
input 	waitrequest;
input 	mem_used_11;
input 	mem_used_12;
input 	waitrequest1;
input 	mem_used_13;
input 	Equal1;
input 	wait_latency_counter_1;
input 	av_readdatavalid;
input 	src_valid;
input 	Equal0;
input 	src_channel_6;
input 	mem;
input 	Equal6;
input 	Equal2;
input 	take_in_data;
input 	saved_grant_11;
input 	Equal5;
input 	saved_grant_12;
input 	src_channel_5;
input 	in_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \read_accepted~2_combout ;
wire \read_accepted~3_combout ;
wire \read_accepted~4_combout ;
wire \read_accepted~5_combout ;
wire \read_accepted~6_combout ;
wire \read_accepted~7_combout ;
wire \read_accepted~8_combout ;
wire \read_accepted~9_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb uav_read(
	.dataa(gnd),
	.datab(gnd),
	.datac(i_read),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read1),
	.cout());
defparam uav_read.lut_mask = 16'h0FFF;
defparam uav_read.sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(rst1),
	.datab(src_valid),
	.datac(wait_latency_counter_1),
	.datad(mem_used_13),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hFEFF;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~1 (
	.dataa(Equal0),
	.datab(src_channel_6),
	.datac(mem),
	.datad(Equal6),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFEFF;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~2 (
	.dataa(Equal1),
	.datab(saved_grant_11),
	.datac(F_pc_5),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(\read_accepted~2_combout ),
	.cout());
defparam \read_accepted~2 .lut_mask = 16'hEFFF;
defparam \read_accepted~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~3 (
	.dataa(saved_grant_12),
	.datab(gnd),
	.datac(waitrequest),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(\read_accepted~3_combout ),
	.cout());
defparam \read_accepted~3 .lut_mask = 16'hAFFF;
defparam \read_accepted~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~4 (
	.dataa(take_in_data),
	.datab(\read_accepted~2_combout ),
	.datac(Equal5),
	.datad(\read_accepted~3_combout ),
	.cin(gnd),
	.combout(\read_accepted~4_combout ),
	.cout());
defparam \read_accepted~4 .lut_mask = 16'hFFFE;
defparam \read_accepted~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~5 (
	.dataa(\read_accepted~1_combout ),
	.datab(\read_accepted~4_combout ),
	.datac(src_channel_5),
	.datad(in_ready),
	.cin(gnd),
	.combout(\read_accepted~5_combout ),
	.cout());
defparam \read_accepted~5 .lut_mask = 16'hFEFF;
defparam \read_accepted~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~6 (
	.dataa(saved_grant_1),
	.datab(F_pc_2),
	.datac(Equal2),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_accepted~6_combout ),
	.cout());
defparam \read_accepted~6 .lut_mask = 16'hFEFF;
defparam \read_accepted~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~7 (
	.dataa(\read_accepted~0_combout ),
	.datab(\read_accepted~5_combout ),
	.datac(\read_accepted~6_combout ),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\read_accepted~7_combout ),
	.cout());
defparam \read_accepted~7 .lut_mask = 16'hFEFF;
defparam \read_accepted~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~8 (
	.dataa(rst1),
	.datab(gnd),
	.datac(gnd),
	.datad(i_read),
	.cin(gnd),
	.combout(\read_accepted~8_combout ),
	.cout());
defparam \read_accepted~8 .lut_mask = 16'hAAFF;
defparam \read_accepted~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~9 (
	.dataa(read_accepted1),
	.datab(\read_accepted~7_combout ),
	.datac(\read_accepted~8_combout ),
	.datad(av_readdatavalid),
	.cin(gnd),
	.combout(\read_accepted~9_combout ),
	.cout());
defparam \read_accepted~9 .lut_mask = 16'hFEFF;
defparam \read_accepted~9 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_agent (
	saved_grant_0,
	WideOr1,
	out_data_buffer_67,
	nonposted_write_endofpacket,
	src_payload_0,
	mem_used_0,
	mem_107_0,
	read_latency_shift_reg_0,
	mem_used_01,
	rp_valid1,
	WideOr0,
	rf_sink_ready,
	out_data_buffer_66,
	nonposted_write_endofpacket1,
	rp_valid2)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_0;
input 	WideOr1;
input 	out_data_buffer_67;
output 	nonposted_write_endofpacket;
input 	src_payload_0;
input 	mem_used_0;
input 	mem_107_0;
input 	read_latency_shift_reg_0;
input 	mem_used_01;
output 	rp_valid1;
input 	WideOr0;
output 	rf_sink_ready;
input 	out_data_buffer_66;
output 	nonposted_write_endofpacket1;
output 	rp_valid2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altera_merlin_burst_uncompressor uncompressor(
	.mem_used_0(mem_used_0),
	.mem_107_0(mem_107_0),
	.rp_valid(rp_valid1),
	.WideOr0(WideOr0),
	.sink_ready(rf_sink_ready));

cycloneive_lcell_comb \nonposted_write_endofpacket~0 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_67),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(nonposted_write_endofpacket),
	.cout());
defparam \nonposted_write_endofpacket~0 .lut_mask = 16'hEEEE;
defparam \nonposted_write_endofpacket~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rp_valid~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(mem_used_01),
	.cin(gnd),
	.combout(rp_valid1),
	.cout());
defparam \rp_valid~0 .lut_mask = 16'h0FFF;
defparam \rp_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nonposted_write_endofpacket~1 (
	.dataa(WideOr1),
	.datab(nonposted_write_endofpacket),
	.datac(src_payload_0),
	.datad(out_data_buffer_66),
	.cin(gnd),
	.combout(nonposted_write_endofpacket1),
	.cout());
defparam \nonposted_write_endofpacket~1 .lut_mask = 16'hFEFF;
defparam \nonposted_write_endofpacket~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb rp_valid(
	.dataa(read_latency_shift_reg_0),
	.datab(mem_used_01),
	.datac(mem_used_0),
	.datad(mem_107_0),
	.cin(gnd),
	.combout(rp_valid2),
	.cout());
defparam rp_valid.lut_mask = 16'hFFFE;
defparam rp_valid.sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_burst_uncompressor (
	mem_used_0,
	mem_107_0,
	rp_valid,
	WideOr0,
	sink_ready)/* synthesis synthesis_greybox=1 */;
input 	mem_used_0;
input 	mem_107_0;
input 	rp_valid;
input 	WideOr0;
output 	sink_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \sink_ready~0 (
	.dataa(mem_used_0),
	.datab(mem_107_0),
	.datac(rp_valid),
	.datad(WideOr0),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hEFFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_agent_1 (
	mem_used_1,
	WideOr1,
	src_data_68,
	m0_read1)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	WideOr1;
input 	src_data_68;
output 	m0_read1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb m0_read(
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(WideOr1),
	.datad(src_data_68),
	.cin(gnd),
	.combout(m0_read1),
	.cout());
defparam m0_read.lut_mask = 16'hAFFF;
defparam m0_read.sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_agent_5 (
	WideOr1,
	mem,
	local_read)/* synthesis synthesis_greybox=1 */;
input 	WideOr1;
input 	mem;
output 	local_read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \local_read~0 (
	.dataa(WideOr1),
	.datab(mem),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(local_read),
	.cout());
defparam \local_read~0 .lut_mask = 16'hEEEE;
defparam \local_read~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_agent_8 (
	mem_used_7,
	saved_grant_0,
	WideOr1,
	out_data_buffer_67,
	src_payload,
	src_payload_0,
	out_data_buffer_66,
	nonposted_write_endofpacket,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	mem_used_7;
input 	saved_grant_0;
input 	WideOr1;
input 	out_data_buffer_67;
input 	src_payload;
input 	src_payload_0;
input 	out_data_buffer_66;
output 	nonposted_write_endofpacket;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \nonposted_write_endofpacket~0 (
	.dataa(WideOr1),
	.datab(src_payload),
	.datac(src_payload_0),
	.datad(out_data_buffer_66),
	.cin(gnd),
	.combout(nonposted_write_endofpacket),
	.cout());
defparam \nonposted_write_endofpacket~0 .lut_mask = 16'hFEFF;
defparam \nonposted_write_endofpacket~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_write~2 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_67),
	.datac(WideOr1),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~2 .lut_mask = 16'hFF7F;
defparam \m0_write~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_agent_9 (
	d_write,
	write_accepted,
	rst1,
	saved_grant_0,
	mem_used_1,
	m0_write,
	wait_latency_counter_1,
	cp_ready)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	rst1;
input 	saved_grant_0;
input 	mem_used_1;
output 	m0_write;
input 	wait_latency_counter_1;
output 	cp_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(write_accepted),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hEFFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cp_ready~0 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(rst1),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(cp_ready),
	.cout());
defparam \cp_ready~0 .lut_mask = 16'hAFFF;
defparam \cp_ready~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator (
	clk,
	reset,
	WideOr1,
	mem_used_1,
	waitrequest_reset_override1,
	read_latency_shift_reg_0,
	src_data_68)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	WideOr1;
input 	mem_used_1;
output 	waitrequest_reset_override1;
output 	read_latency_shift_reg_0;
input 	src_data_68;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas waitrequest_reset_override(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest_reset_override1),
	.prn(vcc));
defparam waitrequest_reset_override.is_wysiwyg = "true";
defparam waitrequest_reset_override.power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(WideOr1),
	.datab(waitrequest_reset_override1),
	.datac(src_data_68),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_1 (
	reset,
	read_latency_shift_reg_0,
	rst1,
	waitrequest,
	m0_read,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	read_latency_shift_reg_0;
input 	rst1;
input 	waitrequest;
input 	m0_read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(gnd),
	.datac(m0_read),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hAFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_2 (
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	d_read,
	read_accepted,
	reset,
	Equal2,
	read_latency_shift_reg_0,
	rst1,
	Equal21,
	av_waitrequest,
	mem_used_1,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	b_full,
	read_0,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_31,
	counter_reg_bit_21,
	counter_reg_bit_01,
	counter_reg_bit_11,
	counter_reg_bit_41,
	counter_reg_bit_51,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_22;
output 	av_readdata_pre_21;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
input 	d_read;
input 	read_accepted;
input 	reset;
input 	Equal2;
output 	read_latency_shift_reg_0;
input 	rst1;
input 	Equal21;
input 	av_waitrequest;
input 	mem_used_1;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
input 	[31:0] av_readdata;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
input 	b_full;
input 	read_0;
input 	counter_reg_bit_3;
input 	counter_reg_bit_0;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	b_full1;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_31;
input 	counter_reg_bit_21;
input 	counter_reg_bit_01;
input 	counter_reg_bit_11;
input 	counter_reg_bit_41;
input 	counter_reg_bit_51;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdata_pre[16]~7_combout ;
wire \av_readdata_pre[16]~8 ;
wire \av_readdata_pre[17]~9_combout ;
wire \av_readdata_pre[17]~10 ;
wire \av_readdata_pre[18]~12 ;
wire \av_readdata_pre[19]~14 ;
wire \av_readdata_pre[20]~16 ;
wire \av_readdata_pre[21]~18 ;
wire \av_readdata_pre[22]~19_combout ;
wire \av_readdata_pre[21]~17_combout ;
wire \av_readdata_pre[20]~15_combout ;
wire \av_readdata_pre[19]~13_combout ;
wire \av_readdata_pre[18]~11_combout ;
wire \read_latency_shift_reg~3_combout ;
wire \av_readdata_pre[13]~21_combout ;


dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(\av_readdata_pre[16]~7_combout ),
	.asdata(counter_reg_bit_01),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(\av_readdata_pre[17]~9_combout ),
	.asdata(counter_reg_bit_11),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(\av_readdata_pre[22]~19_combout ),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(\av_readdata_pre[21]~17_combout ),
	.asdata(counter_reg_bit_51),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(\av_readdata_pre[20]~15_combout ),
	.asdata(counter_reg_bit_41),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(\av_readdata_pre[19]~13_combout ),
	.asdata(counter_reg_bit_31),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(\av_readdata_pre[18]~11_combout ),
	.asdata(counter_reg_bit_21),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(Equal2),
	.datab(Equal21),
	.datac(av_waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

cycloneive_lcell_comb \av_readdata_pre[16]~7 (
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\av_readdata_pre[16]~7_combout ),
	.cout(\av_readdata_pre[16]~8 ));
defparam \av_readdata_pre[16]~7 .lut_mask = 16'hAA55;
defparam \av_readdata_pre[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[17]~9 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[16]~8 ),
	.combout(\av_readdata_pre[17]~9_combout ),
	.cout(\av_readdata_pre[17]~10 ));
defparam \av_readdata_pre[17]~9 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[17]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[18]~11 (
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[17]~10 ),
	.combout(\av_readdata_pre[18]~11_combout ),
	.cout(\av_readdata_pre[18]~12 ));
defparam \av_readdata_pre[18]~11 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[18]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[19]~13 (
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[18]~12 ),
	.combout(\av_readdata_pre[19]~13_combout ),
	.cout(\av_readdata_pre[19]~14 ));
defparam \av_readdata_pre[19]~13 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[19]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[20]~15 (
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[19]~14 ),
	.combout(\av_readdata_pre[20]~15_combout ),
	.cout(\av_readdata_pre[20]~16 ));
defparam \av_readdata_pre[20]~15 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[20]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[21]~17 (
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[20]~16 ),
	.combout(\av_readdata_pre[21]~17_combout ),
	.cout(\av_readdata_pre[21]~18 ));
defparam \av_readdata_pre[21]~17 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[21]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[22]~19 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\av_readdata_pre[21]~18 ),
	.combout(\av_readdata_pre[22]~19_combout ),
	.cout());
defparam \av_readdata_pre[22]~19 .lut_mask = 16'h5A5A;
defparam \av_readdata_pre[22]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \read_latency_shift_reg~3 (
	.dataa(d_read),
	.datab(read_accepted),
	.datac(rst1),
	.datad(read_latency_shift_reg),
	.cin(gnd),
	.combout(\read_latency_shift_reg~3_combout ),
	.cout());
defparam \read_latency_shift_reg~3 .lut_mask = 16'hFFFB;
defparam \read_latency_shift_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[13]~21 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_readdata_pre[13]~21_combout ),
	.cout());
defparam \av_readdata_pre[13]~21 .lut_mask = 16'h5555;
defparam \av_readdata_pre[13]~21 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_3 (
	cp_valid,
	uav_write,
	reset,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	uav_read,
	read_latency_shift_reg_0,
	rst1,
	wait_latency_counter_01,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	cp_valid;
input 	uav_write;
input 	reset;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	uav_read;
output 	read_latency_shift_reg_0;
input 	rst1;
output 	wait_latency_counter_01;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(wait_latency_counter_0),
	.datab(uav_write),
	.datac(always0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(wait_latency_counter_01),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'h96FF;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(uav_read),
	.datab(always0),
	.datac(rst1),
	.datad(wait_latency_counter_01),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(cp_valid),
	.datab(always0),
	.datac(rst1),
	.datad(wait_latency_counter_01),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.cout());
defparam \wait_latency_counter[0]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[0]~1_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[0]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_4 (
	cp_valid,
	uav_write,
	reset,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	uav_read,
	read_latency_shift_reg_0,
	rst1,
	wait_latency_counter_01,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	cp_valid;
input 	uav_write;
input 	reset;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	uav_read;
output 	read_latency_shift_reg_0;
input 	rst1;
output 	wait_latency_counter_01;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter~3_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(wait_latency_counter_0),
	.datab(uav_write),
	.datac(always0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(wait_latency_counter_01),
	.cout());
defparam \wait_latency_counter[0]~0 .lut_mask = 16'h96FF;
defparam \wait_latency_counter[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(uav_read),
	.datab(always0),
	.datac(rst1),
	.datad(wait_latency_counter_01),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(cp_valid),
	.datab(always0),
	.datac(rst1),
	.datad(wait_latency_counter_01),
	.cin(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.cout());
defparam \wait_latency_counter[0]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[0]~1_combout ),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hAFFA;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(wait_latency_counter_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\wait_latency_counter[0]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFF55;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_5 (
	av_readdata,
	reset,
	read_latency_shift_reg_0,
	rst1,
	waitrequest,
	mem_used_1,
	local_read,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_21,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_31,
	av_readdata_pre_30,
	av_readdata_pre_29,
	av_readdata_pre_28,
	av_readdata_pre_27,
	av_readdata_pre_26,
	av_readdata_pre_25,
	av_readdata_pre_10,
	av_readdata_pre_24,
	av_readdata_pre_9,
	av_readdata_pre_23,
	av_readdata_pre_8,
	av_readdata_pre_22,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_20,
	av_readdata_pre_19,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
output 	read_latency_shift_reg_0;
input 	rst1;
input 	waitrequest;
input 	mem_used_1;
input 	local_read;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_11;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	av_readdata_pre_5;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_21;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_31;
output 	av_readdata_pre_30;
output 	av_readdata_pre_29;
output 	av_readdata_pre_28;
output 	av_readdata_pre_27;
output 	av_readdata_pre_26;
output 	av_readdata_pre_25;
output 	av_readdata_pre_10;
output 	av_readdata_pre_24;
output 	av_readdata_pre_9;
output 	av_readdata_pre_23;
output 	av_readdata_pre_8;
output 	av_readdata_pre_22;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(local_read),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_6 (
	reset,
	read_latency_shift_reg_0,
	rst1,
	mem_used_1,
	WideOr1,
	mem,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	read_latency_shift_reg_0;
input 	rst1;
input 	mem_used_1;
input 	WideOr1;
input 	mem;
output 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(mem),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_slave_translator_7 (
	reset,
	read_latency_shift_reg_0,
	rst1,
	mem_used_1,
	WideOr1,
	mem,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	read_latency_shift_reg_0;
input 	rst1;
input 	mem_used_1;
input 	WideOr1;
input 	mem;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(mem),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

endmodule

module final_project_soc_altera_merlin_slave_translator_9 (
	reset,
	read_latency_shift_reg_0,
	rst1,
	mem_used_1,
	WideOr1,
	m0_write,
	wait_latency_counter_1,
	src_data_68,
	read_latency_shift_reg,
	src_payload,
	av_readdata_pre_30,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	read_latency_shift_reg_0;
input 	rst1;
input 	mem_used_1;
input 	WideOr1;
input 	m0_write;
output 	wait_latency_counter_1;
input 	src_data_68;
output 	read_latency_shift_reg;
input 	src_payload;
output 	av_readdata_pre_30;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;
wire \wait_latency_counter[1]~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \wait_latency_counter[0]~q ;
wire \Add0~0_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter[1]~q ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(WideOr1),
	.datac(m0_write),
	.datad(\wait_latency_counter[1]~q ),
	.cin(gnd),
	.combout(wait_latency_counter_1),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'h96FF;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(WideOr1),
	.datac(wait_latency_counter_1),
	.datad(src_data_68),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(read_latency_shift_reg),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hAAFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(rst1),
	.datab(src_payload),
	.datac(src_data_68),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\wait_latency_counter[1]~1_combout ),
	.cout());
defparam \wait_latency_counter[1]~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(\wait_latency_counter[0]~q ),
	.datab(wait_latency_counter_1),
	.datac(WideOr1),
	.datad(\wait_latency_counter[1]~1_combout ),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wait_latency_counter[1]~q ),
	.datad(\wait_latency_counter[0]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~3 (
	.dataa(WideOr1),
	.datab(\Add0~0_combout ),
	.datac(\wait_latency_counter[1]~1_combout ),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.cout());
defparam \wait_latency_counter~3 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter~3 .sum_lutc_input = "datac";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[1]~q ),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_demux (
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	saved_grant_0,
	uav_write,
	mem_used_1,
	Equal0,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	always01,
	wait_latency_counter_11,
	wait_latency_counter_01,
	rst1,
	always1,
	Equal8,
	src_channel_6,
	Equal01,
	src_channel_9,
	in_ready,
	WideOr0,
	read_latency_shift_reg,
	Equal3,
	take_in_data,
	saved_grant_01,
	waitrequest,
	mem_used_11,
	Equal1,
	saved_grant_02,
	mem_used_12,
	saved_grant_03,
	mem_used_13,
	WideOr01,
	saved_grant_04,
	waitrequest1,
	cp_ready,
	WideOr02,
	WideOr03)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_28;
input 	W_alu_result_27;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	saved_grant_0;
input 	uav_write;
input 	mem_used_1;
input 	Equal0;
input 	always0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	always01;
input 	wait_latency_counter_11;
input 	wait_latency_counter_01;
input 	rst1;
input 	always1;
input 	Equal8;
input 	src_channel_6;
input 	Equal01;
input 	src_channel_9;
input 	in_ready;
output 	WideOr0;
input 	read_latency_shift_reg;
input 	Equal3;
input 	take_in_data;
input 	saved_grant_01;
input 	waitrequest;
input 	mem_used_11;
input 	Equal1;
input 	saved_grant_02;
input 	mem_used_12;
input 	saved_grant_03;
input 	mem_used_13;
output 	WideOr01;
input 	saved_grant_04;
input 	waitrequest1;
input 	cp_ready;
output 	WideOr02;
output 	WideOr03;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \WideOr0~3_combout ;
wire \WideOr0~4_combout ;
wire \WideOr0~5_combout ;
wire \WideOr0~6_combout ;
wire \WideOr0~7_combout ;
wire \WideOr0~12_combout ;
wire \WideOr0~8_combout ;
wire \sink_ready~1_combout ;
wire \sink_ready~2_combout ;


cycloneive_lcell_comb \WideOr0~2 (
	.dataa(src_channel_6),
	.datab(Equal01),
	.datac(src_channel_9),
	.datad(in_ready),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'h7FFF;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~9 (
	.dataa(\WideOr0~3_combout ),
	.datab(rst1),
	.datac(\WideOr0~4_combout ),
	.datad(\WideOr0~8_combout ),
	.cin(gnd),
	.combout(WideOr01),
	.cout());
defparam \WideOr0~9 .lut_mask = 16'hFFFE;
defparam \WideOr0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~10 (
	.dataa(\sink_ready~1_combout ),
	.datab(\sink_ready~2_combout ),
	.datac(waitrequest1),
	.datad(cp_ready),
	.cin(gnd),
	.combout(WideOr02),
	.cout());
defparam \WideOr0~10 .lut_mask = 16'hEFFF;
defparam \WideOr0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~11 (
	.dataa(W_alu_result_28),
	.datab(src_channel_6),
	.datac(Equal01),
	.datad(W_alu_result_27),
	.cin(gnd),
	.combout(WideOr03),
	.cout());
defparam \WideOr0~11 .lut_mask = 16'hBFFF;
defparam \WideOr0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~0 (
	.dataa(Equal8),
	.datab(saved_grant_01),
	.datac(waitrequest),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(\sink_ready~0_combout ),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hEFFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~3 (
	.dataa(WideOr0),
	.datab(read_latency_shift_reg),
	.datac(take_in_data),
	.datad(\sink_ready~0_combout ),
	.cin(gnd),
	.combout(\WideOr0~3_combout ),
	.cout());
defparam \WideOr0~3 .lut_mask = 16'hFFFE;
defparam \WideOr0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~4 (
	.dataa(Equal0),
	.datab(Equal1),
	.datac(saved_grant_02),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(\WideOr0~4_combout ),
	.cout());
defparam \WideOr0~4 .lut_mask = 16'hFEFF;
defparam \WideOr0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~5 (
	.dataa(uav_write),
	.datab(always01),
	.datac(wait_latency_counter_01),
	.datad(wait_latency_counter_11),
	.cin(gnd),
	.combout(\WideOr0~5_combout ),
	.cout());
defparam \WideOr0~5 .lut_mask = 16'hDEFF;
defparam \WideOr0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~6 (
	.dataa(always0),
	.datab(uav_write),
	.datac(wait_latency_counter_0),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\WideOr0~6_combout ),
	.cout());
defparam \WideOr0~6 .lut_mask = 16'hBEFF;
defparam \WideOr0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~7 (
	.dataa(W_alu_result_27),
	.datab(W_alu_result_28),
	.datac(saved_grant_03),
	.datad(mem_used_13),
	.cin(gnd),
	.combout(\WideOr0~7_combout ),
	.cout());
defparam \WideOr0~7 .lut_mask = 16'hFBFF;
defparam \WideOr0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~12 (
	.dataa(Equal0),
	.datab(W_alu_result_7),
	.datac(W_alu_result_5),
	.datad(\WideOr0~7_combout ),
	.cin(gnd),
	.combout(\WideOr0~12_combout ),
	.cout());
defparam \WideOr0~12 .lut_mask = 16'hFFBF;
defparam \WideOr0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~8 (
	.dataa(src_channel_6),
	.datab(\WideOr0~5_combout ),
	.datac(\WideOr0~6_combout ),
	.datad(\WideOr0~12_combout ),
	.cin(gnd),
	.combout(\WideOr0~8_combout ),
	.cout());
defparam \WideOr0~8 .lut_mask = 16'hFFFD;
defparam \WideOr0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~1 (
	.dataa(saved_grant_0),
	.datab(W_alu_result_4),
	.datac(Equal3),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\sink_ready~1_combout ),
	.cout());
defparam \sink_ready~1 .lut_mask = 16'hFEFF;
defparam \sink_ready~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~2 (
	.dataa(W_alu_result_7),
	.datab(Equal0),
	.datac(saved_grant_04),
	.datad(always1),
	.cin(gnd),
	.combout(\sink_ready~2_combout ),
	.cout());
defparam \sink_ready~2 .lut_mask = 16'hFFFE;
defparam \sink_ready~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_demux_001 (
	Equal5,
	F_pc_10,
	Equal0,
	F_pc_5,
	Equal01,
	i_read,
	read_accepted,
	uav_read,
	F_pc_2,
	F_pc_4,
	F_pc_9,
	src1_valid,
	Equal1,
	Equal02,
	src_channel_6,
	Equal6,
	src3_valid,
	src6_valid,
	src4_valid)/* synthesis synthesis_greybox=1 */;
input 	Equal5;
input 	F_pc_10;
input 	Equal0;
input 	F_pc_5;
input 	Equal01;
input 	i_read;
input 	read_accepted;
input 	uav_read;
input 	F_pc_2;
input 	F_pc_4;
input 	F_pc_9;
output 	src1_valid;
input 	Equal1;
input 	Equal02;
input 	src_channel_6;
input 	Equal6;
output 	src3_valid;
output 	src6_valid;
output 	src4_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src1_valid~0_combout ;


cycloneive_lcell_comb \src1_valid~1 (
	.dataa(Equal5),
	.datab(Equal0),
	.datac(Equal01),
	.datad(\src1_valid~0_combout ),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~1 .lut_mask = 16'hFFFE;
defparam \src1_valid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src3_valid~0 (
	.dataa(uav_read),
	.datab(Equal5),
	.datac(F_pc_10),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(src3_valid),
	.cout());
defparam \src3_valid~0 .lut_mask = 16'hFEFF;
defparam \src3_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src6_valid~0 (
	.dataa(uav_read),
	.datab(Equal02),
	.datac(src_channel_6),
	.datad(Equal6),
	.cin(gnd),
	.combout(src6_valid),
	.cout());
defparam \src6_valid~0 .lut_mask = 16'hFEFF;
defparam \src6_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src4_valid~2 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(Equal1),
	.datad(F_pc_5),
	.cin(gnd),
	.combout(src4_valid),
	.cout());
defparam \src4_valid~2 .lut_mask = 16'hF7FF;
defparam \src4_valid~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(uav_read),
	.datab(F_pc_2),
	.datac(F_pc_4),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(\src1_valid~0_combout ),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFF;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux (
	clk_0,
	altera_reset_synchronizer_int_chain_out,
	saved_grant_0,
	out_data_buffer_3,
	saved_grant_1,
	out_data_buffer_38,
	out_data_buffer_381,
	src_data_38,
	out_data_buffer_39,
	out_data_buffer_391,
	src_data_39,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	WideOr11,
	mem_used_1,
	last_cycle,
	out_data_buffer_31,
	src_payload,
	waitrequest_reset_override,
	out_data_buffer_107,
	out_data_buffer_1071,
	src_payload_0,
	out_data_buffer_68,
	out_data_buffer_681,
	src_data_68,
	out_data_buffer_30,
	src_payload1,
	out_data_buffer_29,
	src_payload2,
	out_data_buffer_28,
	src_payload3,
	out_data_buffer_0,
	out_data_buffer_1,
	out_data_buffer_2,
	out_data_buffer_27,
	src_payload4,
	out_data_buffer_26,
	src_payload5,
	out_data_buffer_25,
	src_payload6,
	out_data_buffer_24,
	src_payload7,
	out_data_buffer_23,
	src_payload8,
	out_data_buffer_22,
	src_payload9,
	out_data_buffer_21,
	src_payload10,
	out_data_buffer_20,
	src_payload11,
	out_data_buffer_19,
	src_payload12,
	out_data_buffer_18,
	src_payload13,
	out_data_buffer_17,
	src_payload14,
	out_data_buffer_16,
	src_payload15,
	out_data_buffer_15,
	src_payload16,
	out_data_buffer_14,
	src_payload17,
	out_data_buffer_13,
	src_payload18,
	out_data_buffer_12,
	src_payload19,
	out_data_buffer_11,
	src_payload20,
	out_data_buffer_10,
	src_payload21,
	out_data_buffer_9,
	src_payload22,
	out_data_buffer_8,
	src_payload23,
	out_data_buffer_7,
	src_payload24,
	out_data_buffer_6,
	src_payload25,
	out_data_buffer_5,
	src_payload26,
	out_data_buffer_4,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31)/* synthesis synthesis_greybox=1 */;
input 	clk_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	saved_grant_0;
input 	out_data_buffer_3;
output 	saved_grant_1;
input 	out_data_buffer_38;
input 	out_data_buffer_381;
output 	src_data_38;
input 	out_data_buffer_39;
input 	out_data_buffer_391;
output 	src_data_39;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
output 	WideOr11;
input 	mem_used_1;
output 	last_cycle;
input 	out_data_buffer_31;
output 	src_payload;
input 	waitrequest_reset_override;
input 	out_data_buffer_107;
input 	out_data_buffer_1071;
output 	src_payload_0;
input 	out_data_buffer_68;
input 	out_data_buffer_681;
output 	src_data_68;
input 	out_data_buffer_30;
output 	src_payload1;
input 	out_data_buffer_29;
output 	src_payload2;
input 	out_data_buffer_28;
output 	src_payload3;
input 	out_data_buffer_0;
input 	out_data_buffer_1;
input 	out_data_buffer_2;
input 	out_data_buffer_27;
output 	src_payload4;
input 	out_data_buffer_26;
output 	src_payload5;
input 	out_data_buffer_25;
output 	src_payload6;
input 	out_data_buffer_24;
output 	src_payload7;
input 	out_data_buffer_23;
output 	src_payload8;
input 	out_data_buffer_22;
output 	src_payload9;
input 	out_data_buffer_21;
output 	src_payload10;
input 	out_data_buffer_20;
output 	src_payload11;
input 	out_data_buffer_19;
output 	src_payload12;
input 	out_data_buffer_18;
output 	src_payload13;
input 	out_data_buffer_17;
output 	src_payload14;
input 	out_data_buffer_16;
output 	src_payload15;
input 	out_data_buffer_15;
output 	src_payload16;
input 	out_data_buffer_14;
output 	src_payload17;
input 	out_data_buffer_13;
output 	src_payload18;
input 	out_data_buffer_12;
output 	src_payload19;
input 	out_data_buffer_11;
output 	src_payload20;
input 	out_data_buffer_10;
output 	src_payload21;
input 	out_data_buffer_9;
output 	src_payload22;
input 	out_data_buffer_8;
output 	src_payload23;
input 	out_data_buffer_7;
output 	src_payload24;
input 	out_data_buffer_6;
output 	src_payload25;
input 	out_data_buffer_5;
output 	src_payload26;
input 	out_data_buffer_4;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \last_cycle~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


final_project_soc_altera_merlin_arbitrator_6 arb(
	.clk(clk_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid1),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.grant_1(\arb|grant[1]~1_combout ));

dffeas \saved_grant[0] (
	.clk(clk_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb \src_data[38] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_38),
	.datad(out_data_buffer_381),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_39),
	.datad(out_data_buffer_391),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'h7FFF;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_valid),
	.datad(out_valid1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \last_cycle~0 (
	.dataa(WideOr11),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(last_cycle),
	.cout());
defparam \last_cycle~0 .lut_mask = 16'hAAFF;
defparam \last_cycle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_107),
	.datad(out_data_buffer_1071),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0] .lut_mask = 16'hFFFE;
defparam \src_payload[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[68] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_68),
	.datad(out_data_buffer_681),
	.cin(gnd),
	.combout(src_data_68),
	.cout());
defparam \src_data[68] .lut_mask = 16'hFFFE;
defparam \src_data[68] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \last_cycle~1 (
	.dataa(WideOr11),
	.datab(waitrequest_reset_override),
	.datac(src_payload_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\last_cycle~1_combout ),
	.cout());
defparam \last_cycle~1 .lut_mask = 16'hFEFF;
defparam \last_cycle~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(\last_cycle~1_combout ),
	.datab(gnd),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hAFFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_1 (
	W_alu_result_4,
	W_alu_result_11,
	W_alu_result_2,
	W_alu_result_3,
	saved_grant_1,
	cp_valid,
	Equal8,
	Equal3,
	Equal0,
	src_valid,
	uav_read,
	src1_valid,
	saved_grant_0,
	mem_used_1,
	internal_reset,
	d_byteenable_0,
	src_data_32,
	F_pc_0,
	src_data_38,
	F_pc_1,
	src_data_39,
	r_sync_rst,
	d_writedata_16,
	d_writedata_17,
	WideOr11,
	uav_read1,
	src_data_68,
	waitrequest,
	Equal2,
	s_serial_transferSTATE_1_PRE_WRITE,
	src_payload,
	src_payload1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_11;
input 	W_alu_result_2;
input 	W_alu_result_3;
output 	saved_grant_1;
input 	cp_valid;
input 	Equal8;
input 	Equal3;
input 	Equal0;
output 	src_valid;
input 	uav_read;
input 	src1_valid;
output 	saved_grant_0;
input 	mem_used_1;
input 	internal_reset;
input 	d_byteenable_0;
output 	src_data_32;
input 	F_pc_0;
output 	src_data_38;
input 	F_pc_1;
output 	src_data_39;
input 	r_sync_rst;
input 	d_writedata_16;
input 	d_writedata_17;
output 	WideOr11;
input 	uav_read1;
output 	src_data_68;
input 	waitrequest;
input 	Equal2;
input 	s_serial_transferSTATE_1_PRE_WRITE;
output 	src_payload;
output 	src_payload1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \update_grant~1_combout ;
wire \update_grant~2_combout ;
wire \src_valid~0_combout ;


final_project_soc_altera_merlin_arbitrator arb(
	.src_valid(src_valid),
	.src1_valid(src1_valid),
	.reset(r_sync_rst),
	.grant_1(\arb|grant[1]~0_combout ),
	.update_grant(\update_grant~2_combout ),
	.grant_0(\arb|grant[0]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~2_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb \src_valid~1 (
	.dataa(cp_valid),
	.datab(Equal8),
	.datac(Equal3),
	.datad(\src_valid~0_combout ),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~1 .lut_mask = 16'hFFFE;
defparam \src_valid~1 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~2_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cycloneive_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(W_alu_result_2),
	.datad(F_pc_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(W_alu_result_3),
	.datad(F_pc_1),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(src_valid),
	.datad(src1_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[68] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(uav_read1),
	.datad(uav_read),
	.cin(gnd),
	.combout(src_data_68),
	.cout());
defparam \src_data[68] .lut_mask = 16'hFFFE;
defparam \src_data[68] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(mem_used_1),
	.datab(saved_grant_1),
	.datac(saved_grant_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFDFD;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(internal_reset),
	.datab(Equal2),
	.datac(s_serial_transferSTATE_1_PRE_WRITE),
	.datad(\update_grant~0_combout ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'hFFF7;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~2 (
	.dataa(waitrequest),
	.datab(WideOr11),
	.datac(\packet_in_progress~q ),
	.datad(\update_grant~1_combout ),
	.cin(gnd),
	.combout(\update_grant~2_combout ),
	.cout());
defparam \update_grant~2 .lut_mask = 16'hDF1F;
defparam \update_grant~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(W_alu_result_4),
	.datab(Equal0),
	.datac(W_alu_result_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hEFEF;
defparam \src_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_arbitrator (
	src_valid,
	src1_valid,
	reset,
	grant_1,
	update_grant,
	grant_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	src_valid;
input 	src1_valid;
input 	reset;
output 	grant_1;
input 	update_grant;
output 	grant_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[1]~0 (
	.dataa(src1_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~0 .lut_mask = 16'hEFFF;
defparam \grant[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[0]~1 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src1_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~1 .lut_mask = 16'hEFFF;
defparam \grant[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src1_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_2 (
	W_alu_result_7,
	W_alu_result_2,
	d_write,
	write_accepted,
	F_pc_5,
	i_read,
	read_accepted,
	uav_read,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	Equal0,
	uav_read1,
	rst1,
	always1,
	saved_grant_0,
	mem_used_1,
	Equal1,
	saved_grant_1,
	WideOr11,
	wait_latency_counter_1,
	always11,
	src_valid,
	src_data_68,
	always12,
	src_payload,
	src_data_38,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_2;
input 	d_write;
input 	write_accepted;
input 	F_pc_5;
input 	i_read;
input 	read_accepted;
input 	uav_read;
input 	F_pc_0;
input 	F_pc_1;
input 	r_sync_rst;
input 	Equal0;
input 	uav_read1;
input 	rst1;
input 	always1;
output 	saved_grant_0;
input 	mem_used_1;
input 	Equal1;
output 	saved_grant_1;
output 	WideOr11;
input 	wait_latency_counter_1;
input 	always11;
output 	src_valid;
output 	src_data_68;
input 	always12;
output 	src_payload;
output 	src_data_38;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~2_combout ;
wire \arb|grant[1]~4_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \update_grant~1_combout ;
wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;


final_project_soc_altera_merlin_arbitrator_1 arb(
	.i_read(i_read),
	.read_accepted(read_accepted),
	.reset(r_sync_rst),
	.always1(always11),
	.always11(always12),
	.grant_0(\arb|grant[0]~2_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~4_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(Equal0),
	.datab(Equal1),
	.datac(\WideOr1~0_combout ),
	.datad(\WideOr1~1_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(saved_grant_1),
	.datab(always11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hEEEE;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[68] (
	.dataa(uav_read),
	.datab(uav_read1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_68),
	.cout());
defparam \src_data[68] .lut_mask = 16'hFFFE;
defparam \src_data[68] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(d_write),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(mem_used_1),
	.datab(rst1),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFFFD;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(WideOr11),
	.datab(\packet_in_progress~q ),
	.datac(wait_latency_counter_1),
	.datad(\update_grant~0_combout ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'hF7B3;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(saved_grant_1),
	.datab(uav_read),
	.datac(F_pc_5),
	.datad(F_pc_1),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~1 (
	.dataa(saved_grant_0),
	.datab(W_alu_result_7),
	.datac(always1),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr1~1_combout ),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'hFEFE;
defparam \WideOr1~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_arbitrator_1 (
	i_read,
	read_accepted,
	reset,
	always1,
	always11,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	i_read;
input 	read_accepted;
input 	reset;
input 	always1;
input 	always11;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;
wire \grant[1]~3_combout ;


cycloneive_lcell_comb \grant[0]~2 (
	.dataa(always11),
	.datab(\top_priority_reg[1]~q ),
	.datac(always1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~2 .lut_mask = 16'hEFFF;
defparam \grant[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~4 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(always1),
	.datad(\grant[1]~3_combout ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~4 .lut_mask = 16'hFFF7;
defparam \grant[1]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(always11),
	.datac(always1),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

cycloneive_lcell_comb \grant[1]~3 (
	.dataa(\top_priority_reg[1]~q ),
	.datab(gnd),
	.datac(always11),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(\grant[1]~3_combout ),
	.cout());
defparam \grant[1]~3 .lut_mask = 16'hAFFF;
defparam \grant[1]~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_3 (
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_11,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	cp_valid,
	Equal8,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_3,
	F_pc_2,
	F_pc_4,
	d_writedata_0,
	d_byteenable_0,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_1,
	src3_valid,
	WideOr11,
	hbreak_enabled,
	d_byteenable_2,
	src_data_46,
	d_byteenable_1,
	d_byteenable_3,
	d_writedata_21,
	d_writedata_18,
	d_writedata_23,
	d_writedata_22,
	d_writedata_20,
	d_writedata_19,
	src_payload,
	src_payload1,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_33,
	src_payload7,
	src_payload8,
	src_data_34,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_35,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_12;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_11;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_31;
input 	d_writedata_30;
input 	d_writedata_29;
input 	d_writedata_28;
input 	d_writedata_27;
input 	d_writedata_26;
input 	d_writedata_25;
input 	d_writedata_24;
input 	cp_valid;
input 	Equal8;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_3;
input 	F_pc_2;
input 	F_pc_4;
input 	d_writedata_0;
input 	d_byteenable_0;
input 	F_pc_0;
input 	F_pc_1;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
output 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
output 	saved_grant_1;
input 	src3_valid;
output 	WideOr11;
input 	hbreak_enabled;
input 	d_byteenable_2;
output 	src_data_46;
input 	d_byteenable_1;
input 	d_byteenable_3;
input 	d_writedata_21;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_22;
input 	d_writedata_20;
input 	d_writedata_19;
output 	src_payload;
output 	src_payload1;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_data_33;
output 	src_payload7;
output 	src_payload8;
output 	src_data_34;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_data_35;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~0_combout ;


final_project_soc_altera_merlin_arbitrator_2 arb(
	.reset(r_sync_rst),
	.src_valid(\src_valid~0_combout ),
	.src3_valid(src3_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_valid~0_combout ),
	.datad(src3_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(F_pc_8),
	.datab(W_alu_result_10),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(F_pc_2),
	.datab(W_alu_result_4),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(F_pc_3),
	.datab(W_alu_result_5),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(F_pc_4),
	.datab(W_alu_result_6),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(F_pc_5),
	.datab(W_alu_result_7),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(F_pc_6),
	.datab(W_alu_result_8),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(F_pc_7),
	.datab(W_alu_result_9),
	.datac(saved_grant_0),
	.datad(saved_grant_1),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(d_byteenable_0),
	.datac(saved_grant_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(d_writedata_11),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(d_writedata_13),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(d_writedata_16),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(d_writedata_12),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(d_writedata_14),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(d_writedata_15),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(d_writedata_17),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(d_writedata_10),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(d_writedata_9),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(d_writedata_8),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEFFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(cp_valid),
	.datab(Equal8),
	.datac(W_alu_result_12),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hFEFF;
defparam \src_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_arbitrator_2 (
	reset,
	src_valid,
	src3_valid,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src_valid;
input 	src3_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src3_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src3_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src3_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_4 (
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	cp_valid,
	F_pc_5,
	i_read,
	read_accepted,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	Equal0,
	rst1,
	saved_grant_0,
	mem_used_1,
	Equal1,
	saved_grant_1,
	WideOr11,
	src_data_38,
	src_data_39,
	src4_valid,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	cp_valid;
input 	F_pc_5;
input 	i_read;
input 	read_accepted;
input 	F_pc_0;
input 	F_pc_1;
input 	r_sync_rst;
input 	Equal0;
input 	rst1;
output 	saved_grant_0;
input 	mem_used_1;
input 	Equal1;
output 	saved_grant_1;
output 	WideOr11;
output 	src_data_38;
output 	src_data_39;
input 	src4_valid;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_valid~0_combout ;
wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \WideOr1~2_combout ;
wire \WideOr1~3_combout ;


final_project_soc_altera_merlin_arbitrator_3 arb(
	.reset(r_sync_rst),
	.src_valid(\src_valid~0_combout ),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.src4_valid(src4_valid),
	.clk(clk_clk));

cycloneive_lcell_comb \src_valid~0 (
	.dataa(cp_valid),
	.datab(W_alu_result_5),
	.datac(Equal0),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hFEFF;
defparam \src_valid~0 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(Equal0),
	.datab(Equal1),
	.datac(\WideOr1~2_combout ),
	.datad(\WideOr1~3_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(rst1),
	.datab(saved_grant_1),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFEFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~2 (
	.dataa(saved_grant_0),
	.datab(cp_valid),
	.datac(W_alu_result_5),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(\WideOr1~2_combout ),
	.cout());
defparam \WideOr1~2 .lut_mask = 16'hFEFF;
defparam \WideOr1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~3 (
	.dataa(i_read),
	.datab(read_accepted),
	.datac(saved_grant_1),
	.datad(F_pc_5),
	.cin(gnd),
	.combout(\WideOr1~3_combout ),
	.cout());
defparam \WideOr1~3 .lut_mask = 16'hF7FF;
defparam \WideOr1~3 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_arbitrator_3 (
	reset,
	src_valid,
	grant_0,
	update_grant,
	grant_1,
	src4_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	src4_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src4_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src4_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src4_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_5 (
	wire_pll7_clk_0,
	entries_1,
	entries_0,
	altera_reset_synchronizer_int_chain_out,
	mem_used_7,
	last_cycle,
	saved_grant_0,
	saved_grant_1,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	WideOr11,
	out_data_buffer_67,
	src_payload,
	out_data_buffer_68,
	out_data_buffer_681,
	src_data_68,
	out_data_buffer_48,
	out_data_buffer_481,
	src_data_48,
	out_data_buffer_62,
	out_data_buffer_621,
	src_data_62,
	out_data_buffer_49,
	out_data_buffer_491,
	src_data_49,
	out_data_buffer_51,
	out_data_buffer_511,
	src_data_51,
	out_data_buffer_50,
	out_data_buffer_501,
	src_data_50,
	out_data_buffer_53,
	out_data_buffer_531,
	src_data_53,
	out_data_buffer_52,
	out_data_buffer_521,
	src_data_52,
	out_data_buffer_55,
	out_data_buffer_551,
	src_data_55,
	out_data_buffer_54,
	out_data_buffer_541,
	src_data_54,
	out_data_buffer_57,
	out_data_buffer_571,
	src_data_57,
	out_data_buffer_56,
	out_data_buffer_561,
	src_data_56,
	out_data_buffer_59,
	out_data_buffer_591,
	src_data_59,
	out_data_buffer_58,
	out_data_buffer_581,
	src_data_58,
	out_data_buffer_61,
	out_data_buffer_611,
	src_data_61,
	out_data_buffer_60,
	out_data_buffer_601,
	src_data_60,
	out_data_buffer_38,
	out_data_buffer_381,
	src_data_38,
	out_data_buffer_39,
	out_data_buffer_391,
	src_data_39,
	out_data_buffer_40,
	out_data_buffer_401,
	src_data_40,
	out_data_buffer_41,
	out_data_buffer_411,
	src_data_41,
	out_data_buffer_42,
	out_data_buffer_421,
	src_data_42,
	out_data_buffer_43,
	out_data_buffer_431,
	src_data_43,
	out_data_buffer_44,
	out_data_buffer_441,
	src_data_44,
	out_data_buffer_45,
	out_data_buffer_451,
	src_data_45,
	out_data_buffer_46,
	out_data_buffer_461,
	src_data_46,
	out_data_buffer_47,
	out_data_buffer_471,
	src_data_47,
	out_data_buffer_107,
	out_data_buffer_1071,
	src_payload_0,
	out_data_buffer_0,
	src_payload1,
	out_data_buffer_1,
	src_payload2,
	out_data_buffer_2,
	src_payload3,
	out_data_buffer_3,
	src_payload4,
	out_data_buffer_4,
	src_payload5,
	out_data_buffer_5,
	src_payload6,
	out_data_buffer_6,
	src_payload7,
	out_data_buffer_7,
	src_payload8,
	out_data_buffer_8,
	src_payload9,
	out_data_buffer_9,
	src_payload10,
	out_data_buffer_10,
	src_payload11,
	out_data_buffer_11,
	src_payload12,
	out_data_buffer_12,
	src_payload13,
	out_data_buffer_13,
	src_payload14,
	out_data_buffer_14,
	src_payload15,
	out_data_buffer_15,
	src_payload16,
	out_data_buffer_16,
	src_payload17,
	out_data_buffer_17,
	src_payload18,
	out_data_buffer_18,
	src_payload19,
	out_data_buffer_19,
	src_payload20,
	out_data_buffer_20,
	src_payload21,
	out_data_buffer_21,
	src_payload22,
	out_data_buffer_22,
	src_payload23,
	out_data_buffer_23,
	src_payload24,
	out_data_buffer_24,
	src_payload25,
	out_data_buffer_25,
	src_payload26,
	out_data_buffer_26,
	src_payload27,
	out_data_buffer_27,
	src_payload28,
	out_data_buffer_28,
	src_payload29,
	out_data_buffer_29,
	src_payload30,
	out_data_buffer_30,
	src_payload31,
	out_data_buffer_31,
	src_payload32)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
input 	entries_1;
input 	entries_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	mem_used_7;
output 	last_cycle;
output 	saved_grant_0;
output 	saved_grant_1;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
output 	WideOr11;
input 	out_data_buffer_67;
output 	src_payload;
input 	out_data_buffer_68;
input 	out_data_buffer_681;
output 	src_data_68;
input 	out_data_buffer_48;
input 	out_data_buffer_481;
output 	src_data_48;
input 	out_data_buffer_62;
input 	out_data_buffer_621;
output 	src_data_62;
input 	out_data_buffer_49;
input 	out_data_buffer_491;
output 	src_data_49;
input 	out_data_buffer_51;
input 	out_data_buffer_511;
output 	src_data_51;
input 	out_data_buffer_50;
input 	out_data_buffer_501;
output 	src_data_50;
input 	out_data_buffer_53;
input 	out_data_buffer_531;
output 	src_data_53;
input 	out_data_buffer_52;
input 	out_data_buffer_521;
output 	src_data_52;
input 	out_data_buffer_55;
input 	out_data_buffer_551;
output 	src_data_55;
input 	out_data_buffer_54;
input 	out_data_buffer_541;
output 	src_data_54;
input 	out_data_buffer_57;
input 	out_data_buffer_571;
output 	src_data_57;
input 	out_data_buffer_56;
input 	out_data_buffer_561;
output 	src_data_56;
input 	out_data_buffer_59;
input 	out_data_buffer_591;
output 	src_data_59;
input 	out_data_buffer_58;
input 	out_data_buffer_581;
output 	src_data_58;
input 	out_data_buffer_61;
input 	out_data_buffer_611;
output 	src_data_61;
input 	out_data_buffer_60;
input 	out_data_buffer_601;
output 	src_data_60;
input 	out_data_buffer_38;
input 	out_data_buffer_381;
output 	src_data_38;
input 	out_data_buffer_39;
input 	out_data_buffer_391;
output 	src_data_39;
input 	out_data_buffer_40;
input 	out_data_buffer_401;
output 	src_data_40;
input 	out_data_buffer_41;
input 	out_data_buffer_411;
output 	src_data_41;
input 	out_data_buffer_42;
input 	out_data_buffer_421;
output 	src_data_42;
input 	out_data_buffer_43;
input 	out_data_buffer_431;
output 	src_data_43;
input 	out_data_buffer_44;
input 	out_data_buffer_441;
output 	src_data_44;
input 	out_data_buffer_45;
input 	out_data_buffer_451;
output 	src_data_45;
input 	out_data_buffer_46;
input 	out_data_buffer_461;
output 	src_data_46;
input 	out_data_buffer_47;
input 	out_data_buffer_471;
output 	src_data_47;
input 	out_data_buffer_107;
input 	out_data_buffer_1071;
output 	src_payload_0;
input 	out_data_buffer_0;
output 	src_payload1;
input 	out_data_buffer_1;
output 	src_payload2;
input 	out_data_buffer_2;
output 	src_payload3;
input 	out_data_buffer_3;
output 	src_payload4;
input 	out_data_buffer_4;
output 	src_payload5;
input 	out_data_buffer_5;
output 	src_payload6;
input 	out_data_buffer_6;
output 	src_payload7;
input 	out_data_buffer_7;
output 	src_payload8;
input 	out_data_buffer_8;
output 	src_payload9;
input 	out_data_buffer_9;
output 	src_payload10;
input 	out_data_buffer_10;
output 	src_payload11;
input 	out_data_buffer_11;
output 	src_payload12;
input 	out_data_buffer_12;
output 	src_payload13;
input 	out_data_buffer_13;
output 	src_payload14;
input 	out_data_buffer_14;
output 	src_payload15;
input 	out_data_buffer_15;
output 	src_payload16;
input 	out_data_buffer_16;
output 	src_payload17;
input 	out_data_buffer_17;
output 	src_payload18;
input 	out_data_buffer_18;
output 	src_payload19;
input 	out_data_buffer_19;
output 	src_payload20;
input 	out_data_buffer_20;
output 	src_payload21;
input 	out_data_buffer_21;
output 	src_payload22;
input 	out_data_buffer_22;
output 	src_payload23;
input 	out_data_buffer_23;
output 	src_payload24;
input 	out_data_buffer_24;
output 	src_payload25;
input 	out_data_buffer_25;
output 	src_payload26;
input 	out_data_buffer_26;
output 	src_payload27;
input 	out_data_buffer_27;
output 	src_payload28;
input 	out_data_buffer_28;
output 	src_payload29;
input 	out_data_buffer_29;
output 	src_payload30;
input 	out_data_buffer_30;
output 	src_payload31;
input 	out_data_buffer_31;
output 	src_payload32;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


final_project_soc_altera_merlin_arbitrator_4 arb(
	.clk(wire_pll7_clk_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid1),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.grant_1(\arb|grant[1]~1_combout ));

cycloneive_lcell_comb \last_cycle~0 (
	.dataa(entries_0),
	.datab(gnd),
	.datac(entries_1),
	.datad(mem_used_7),
	.cin(gnd),
	.combout(last_cycle),
	.cout());
defparam \last_cycle~0 .lut_mask = 16'hAFFF;
defparam \last_cycle~0 .sum_lutc_input = "datac";

dffeas \saved_grant[0] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(wire_pll7_clk_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_valid),
	.datad(out_valid1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_67),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[68] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_68),
	.datad(out_data_buffer_681),
	.cin(gnd),
	.combout(src_data_68),
	.cout());
defparam \src_data[68] .lut_mask = 16'hFFFE;
defparam \src_data[68] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[48] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_48),
	.datad(out_data_buffer_481),
	.cin(gnd),
	.combout(src_data_48),
	.cout());
defparam \src_data[48] .lut_mask = 16'hFFFE;
defparam \src_data[48] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[62] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_62),
	.datad(out_data_buffer_621),
	.cin(gnd),
	.combout(src_data_62),
	.cout());
defparam \src_data[62] .lut_mask = 16'hFFFE;
defparam \src_data[62] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[49] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_49),
	.datad(out_data_buffer_491),
	.cin(gnd),
	.combout(src_data_49),
	.cout());
defparam \src_data[49] .lut_mask = 16'hFFFE;
defparam \src_data[49] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[51] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_51),
	.datad(out_data_buffer_511),
	.cin(gnd),
	.combout(src_data_51),
	.cout());
defparam \src_data[51] .lut_mask = 16'hFFFE;
defparam \src_data[51] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[50] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_50),
	.datad(out_data_buffer_501),
	.cin(gnd),
	.combout(src_data_50),
	.cout());
defparam \src_data[50] .lut_mask = 16'hFFFE;
defparam \src_data[50] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[53] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_53),
	.datad(out_data_buffer_531),
	.cin(gnd),
	.combout(src_data_53),
	.cout());
defparam \src_data[53] .lut_mask = 16'hFFFE;
defparam \src_data[53] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[52] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_52),
	.datad(out_data_buffer_521),
	.cin(gnd),
	.combout(src_data_52),
	.cout());
defparam \src_data[52] .lut_mask = 16'hFFFE;
defparam \src_data[52] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[55] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_55),
	.datad(out_data_buffer_551),
	.cin(gnd),
	.combout(src_data_55),
	.cout());
defparam \src_data[55] .lut_mask = 16'hFFFE;
defparam \src_data[55] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[54] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_54),
	.datad(out_data_buffer_541),
	.cin(gnd),
	.combout(src_data_54),
	.cout());
defparam \src_data[54] .lut_mask = 16'hFFFE;
defparam \src_data[54] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[57] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_57),
	.datad(out_data_buffer_571),
	.cin(gnd),
	.combout(src_data_57),
	.cout());
defparam \src_data[57] .lut_mask = 16'hFFFE;
defparam \src_data[57] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[56] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_56),
	.datad(out_data_buffer_561),
	.cin(gnd),
	.combout(src_data_56),
	.cout());
defparam \src_data[56] .lut_mask = 16'hFFFE;
defparam \src_data[56] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[59] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_59),
	.datad(out_data_buffer_591),
	.cin(gnd),
	.combout(src_data_59),
	.cout());
defparam \src_data[59] .lut_mask = 16'hFFFE;
defparam \src_data[59] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[58] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_58),
	.datad(out_data_buffer_581),
	.cin(gnd),
	.combout(src_data_58),
	.cout());
defparam \src_data[58] .lut_mask = 16'hFFFE;
defparam \src_data[58] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[61] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_61),
	.datad(out_data_buffer_611),
	.cin(gnd),
	.combout(src_data_61),
	.cout());
defparam \src_data[61] .lut_mask = 16'hFFFE;
defparam \src_data[61] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[60] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_60),
	.datad(out_data_buffer_601),
	.cin(gnd),
	.combout(src_data_60),
	.cout());
defparam \src_data[60] .lut_mask = 16'hFFFE;
defparam \src_data[60] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_38),
	.datad(out_data_buffer_381),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_39),
	.datad(out_data_buffer_391),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_40),
	.datad(out_data_buffer_401),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_41),
	.datad(out_data_buffer_411),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_42),
	.datad(out_data_buffer_421),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_43),
	.datad(out_data_buffer_431),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_44),
	.datad(out_data_buffer_441),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_45),
	.datad(out_data_buffer_451),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_46),
	.datad(out_data_buffer_461),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[47] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_47),
	.datad(out_data_buffer_471),
	.cin(gnd),
	.combout(src_data_47),
	.cout());
defparam \src_data[47] .lut_mask = 16'hFFFE;
defparam \src_data[47] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0] (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(out_data_buffer_107),
	.datad(out_data_buffer_1071),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0] .lut_mask = 16'hFFFE;
defparam \src_payload[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(out_data_buffer_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(wire_pll7_clk_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(last_cycle),
	.datab(src_payload_0),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hACFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_arbitrator_4 (
	clk,
	reset,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	grant_0,
	update_grant,
	grant_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
output 	grant_0;
input 	update_grant;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~4_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~5_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(out_valid1),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(out_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~4 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(update_grant),
	.datad(out_valid),
	.cin(gnd),
	.combout(\top_priority_reg[0]~4_combout ),
	.cout());
defparam \top_priority_reg[0]~4 .lut_mask = 16'hFFF6;
defparam \top_priority_reg[0]~4 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~5 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~5_combout ),
	.cout());
defparam \top_priority_reg[0]~5 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~5 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_cmd_mux_6 (
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_2,
	W_alu_result_3,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	cp_valid,
	d_writedata_0,
	d_byteenable_0,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	Equal0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	rst1,
	src_channel_6,
	src_channel_61,
	Equal8,
	Equal2,
	src_channel_9,
	saved_grant_0,
	mem_used_1,
	saved_grant_1,
	src6_valid,
	WideOr11,
	d_byteenable_2,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_32,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	d_byteenable_1,
	d_byteenable_3,
	src_payload5,
	src_data_33,
	src_payload6,
	src_payload7,
	src_data_34,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	d_writedata_21,
	src_payload12,
	d_writedata_18,
	src_payload13,
	src_payload14,
	src_payload15,
	src_data_35,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	d_writedata_23,
	src_payload25,
	src_payload26,
	d_writedata_22,
	src_payload27,
	src_payload28,
	src_payload29,
	d_writedata_20,
	src_payload30,
	d_writedata_19,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_2;
input 	W_alu_result_3;
input 	d_writedata_31;
input 	d_writedata_30;
input 	d_writedata_29;
input 	d_writedata_28;
input 	d_writedata_27;
input 	d_writedata_26;
input 	d_writedata_25;
input 	d_writedata_24;
input 	cp_valid;
input 	d_writedata_0;
input 	d_byteenable_0;
input 	F_pc_0;
input 	F_pc_1;
input 	r_sync_rst;
input 	Equal0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	d_writedata_8;
input 	d_writedata_9;
input 	d_writedata_10;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_17;
input 	rst1;
input 	src_channel_6;
input 	src_channel_61;
input 	Equal8;
input 	Equal2;
input 	src_channel_9;
output 	saved_grant_0;
input 	mem_used_1;
output 	saved_grant_1;
input 	src6_valid;
output 	WideOr11;
input 	d_byteenable_2;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_32;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
input 	d_byteenable_1;
input 	d_byteenable_3;
output 	src_payload5;
output 	src_data_33;
output 	src_payload6;
output 	src_payload7;
output 	src_data_34;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
input 	d_writedata_21;
output 	src_payload12;
input 	d_writedata_18;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_data_35;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
input 	d_writedata_23;
output 	src_payload25;
output 	src_payload26;
input 	d_writedata_22;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
input 	d_writedata_20;
output 	src_payload30;
input 	d_writedata_19;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;
wire \src_valid~0_combout ;
wire \src_valid~1_combout ;
wire \src_valid~2_combout ;


final_project_soc_altera_merlin_arbitrator_5 arb(
	.reset(r_sync_rst),
	.src_valid(\src_valid~2_combout ),
	.src6_valid(src6_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_valid~2_combout ),
	.datad(src6_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(d_byteenable_0),
	.datac(saved_grant_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(d_writedata_11),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(d_writedata_13),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(d_writedata_16),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(d_writedata_12),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(d_writedata_14),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(d_writedata_15),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(d_writedata_17),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(d_writedata_10),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(d_writedata_9),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(d_writedata_8),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(rst1),
	.datab(saved_grant_1),
	.datac(saved_grant_0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hFEFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(cp_valid),
	.datab(src_channel_9),
	.datac(W_alu_result_7),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'hEFFF;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~1 (
	.dataa(src_channel_61),
	.datab(Equal2),
	.datac(\src_valid~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_valid~1_combout ),
	.cout());
defparam \src_valid~1 .lut_mask = 16'hF7F7;
defparam \src_valid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~2 (
	.dataa(src_channel_6),
	.datab(Equal8),
	.datac(Equal0),
	.datad(\src_valid~1_combout ),
	.cin(gnd),
	.combout(\src_valid~2_combout ),
	.cout());
defparam \src_valid~2 .lut_mask = 16'hFFF7;
defparam \src_valid~2 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_merlin_arbitrator_5 (
	reset,
	src_valid,
	src6_valid,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src_valid;
input 	src6_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src6_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src6_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src6_valid),
	.datac(src_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module final_project_soc_altera_merlin_arbitrator_6 (
	clk,
	reset,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	grant_0,
	update_grant,
	grant_1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
output 	grant_0;
input 	update_grant;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~4_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~5_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(out_valid1),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(out_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(out_valid1),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~4 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(update_grant),
	.datad(out_valid),
	.cin(gnd),
	.combout(\top_priority_reg[0]~4_combout ),
	.cout());
defparam \top_priority_reg[0]~4 .lut_mask = 16'hFFF6;
defparam \top_priority_reg[0]~4 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~5 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~5_combout ),
	.cout());
defparam \top_priority_reg[0]~5 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~5 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~4_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_router (
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_11,
	W_alu_result_3,
	d_read,
	read_accepted,
	Equal8,
	Equal3,
	Equal0,
	Equal01,
	Equal2,
	always1,
	src_channel_6,
	src_channel_61,
	Equal81,
	Equal21,
	src_channel_62,
	Equal02,
	src_channel_9,
	Equal22,
	Equal31,
	Equal1,
	always11)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_28;
input 	W_alu_result_27;
input 	W_alu_result_26;
input 	W_alu_result_25;
input 	W_alu_result_24;
input 	W_alu_result_23;
input 	W_alu_result_22;
input 	W_alu_result_21;
input 	W_alu_result_20;
input 	W_alu_result_19;
input 	W_alu_result_18;
input 	W_alu_result_17;
input 	W_alu_result_16;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_6;
input 	W_alu_result_7;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_12;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_11;
input 	W_alu_result_3;
input 	d_read;
input 	read_accepted;
output 	Equal8;
output 	Equal3;
output 	Equal0;
output 	Equal01;
output 	Equal2;
output 	always1;
output 	src_channel_6;
output 	src_channel_61;
output 	Equal81;
output 	Equal21;
output 	src_channel_62;
output 	Equal02;
output 	src_channel_9;
output 	Equal22;
output 	Equal31;
output 	Equal1;
output 	always11;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal8~0_combout ;
wire \Equal8~1_combout ;
wire \Equal8~2_combout ;
wire \Equal8~3_combout ;
wire \Equal0~1_combout ;
wire \Equal2~0_combout ;
wire \src_channel[6]~4_combout ;
wire \src_channel[6]~9_combout ;
wire \Equal2~2_combout ;
wire \always1~1_combout ;


cycloneive_lcell_comb \Equal8~4 (
	.dataa(\Equal8~0_combout ),
	.datab(\Equal8~1_combout ),
	.datac(\Equal8~2_combout ),
	.datad(\Equal8~3_combout ),
	.cin(gnd),
	.combout(Equal8),
	.cout());
defparam \Equal8~4 .lut_mask = 16'hFFFE;
defparam \Equal8~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(W_alu_result_6),
	.datab(gnd),
	.datac(W_alu_result_7),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(Equal3),
	.cout());
defparam \Equal3~0 .lut_mask = 16'hAFFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(W_alu_result_12),
	.datab(W_alu_result_10),
	.datac(W_alu_result_9),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(\Equal0~1_combout ),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(\Equal2~0_combout ),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hFEFF;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(d_read),
	.datab(W_alu_result_5),
	.datac(W_alu_result_3),
	.datad(read_accepted),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~5 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(\Equal0~1_combout ),
	.datad(\src_channel[6]~4_combout ),
	.cin(gnd),
	.combout(src_channel_6),
	.cout());
defparam \src_channel[6]~5 .lut_mask = 16'hFFFE;
defparam \src_channel[6]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~6 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(W_alu_result_11),
	.datad(\src_channel[6]~9_combout ),
	.cin(gnd),
	.combout(src_channel_61),
	.cout());
defparam \src_channel[6]~6 .lut_mask = 16'hFFEF;
defparam \src_channel[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal8~5 (
	.dataa(Equal8),
	.datab(W_alu_result_12),
	.datac(gnd),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(Equal81),
	.cout());
defparam \Equal8~5 .lut_mask = 16'hEEFF;
defparam \Equal8~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~3 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(\Equal2~0_combout ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(Equal21),
	.cout());
defparam \Equal2~3 .lut_mask = 16'hFFFE;
defparam \Equal2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~7 (
	.dataa(src_channel_6),
	.datab(src_channel_61),
	.datac(Equal81),
	.datad(Equal21),
	.cin(gnd),
	.combout(src_channel_62),
	.cout());
defparam \src_channel[6]~7 .lut_mask = 16'hFFFE;
defparam \src_channel[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(Equal01),
	.datab(gnd),
	.datac(W_alu_result_7),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(Equal02),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hAFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[9]~8 (
	.dataa(W_alu_result_27),
	.datab(gnd),
	.datac(gnd),
	.datad(W_alu_result_28),
	.cin(gnd),
	.combout(src_channel_9),
	.cout());
defparam \src_channel[9]~8 .lut_mask = 16'hAAFF;
defparam \src_channel[9]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_6),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(Equal22),
	.cout());
defparam \Equal2~4 .lut_mask = 16'h0FFF;
defparam \Equal2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~1 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(Equal3),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(Equal31),
	.cout());
defparam \Equal3~1 .lut_mask = 16'hFEFF;
defparam \Equal3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(W_alu_result_5),
	.datab(gnd),
	.datac(gnd),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hAAFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~2 (
	.dataa(Equal8),
	.datab(Equal0),
	.datac(\Equal0~1_combout ),
	.datad(\always1~1_combout ),
	.cin(gnd),
	.combout(always11),
	.cout());
defparam \always1~2 .lut_mask = 16'hFFFE;
defparam \always1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal8~0 (
	.dataa(W_alu_result_28),
	.datab(W_alu_result_27),
	.datac(W_alu_result_26),
	.datad(W_alu_result_25),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
defparam \Equal8~0 .lut_mask = 16'h7FFF;
defparam \Equal8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal8~1 (
	.dataa(W_alu_result_24),
	.datab(W_alu_result_23),
	.datac(W_alu_result_22),
	.datad(W_alu_result_21),
	.cin(gnd),
	.combout(\Equal8~1_combout ),
	.cout());
defparam \Equal8~1 .lut_mask = 16'h7FFF;
defparam \Equal8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal8~2 (
	.dataa(W_alu_result_20),
	.datab(W_alu_result_19),
	.datac(W_alu_result_18),
	.datad(W_alu_result_17),
	.cin(gnd),
	.combout(\Equal8~2_combout ),
	.cout());
defparam \Equal8~2 .lut_mask = 16'h7FFF;
defparam \Equal8~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal8~3 (
	.dataa(W_alu_result_16),
	.datab(W_alu_result_15),
	.datac(W_alu_result_14),
	.datad(W_alu_result_13),
	.cin(gnd),
	.combout(\Equal8~3_combout ),
	.cout());
defparam \Equal8~3 .lut_mask = 16'h7FFF;
defparam \Equal8~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_4),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h0FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_5),
	.datac(gnd),
	.datad(W_alu_result_7),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEEFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~4 (
	.dataa(always1),
	.datab(W_alu_result_7),
	.datac(W_alu_result_5),
	.datad(W_alu_result_11),
	.cin(gnd),
	.combout(\src_channel[6]~4_combout ),
	.cout());
defparam \src_channel[6]~4 .lut_mask = 16'hBEFF;
defparam \src_channel[6]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~9 (
	.dataa(W_alu_result_4),
	.datab(W_alu_result_5),
	.datac(W_alu_result_7),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\src_channel[6]~9_combout ),
	.cout());
defparam \src_channel[6]~9 .lut_mask = 16'hFFBF;
defparam \src_channel[6]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~2 (
	.dataa(W_alu_result_6),
	.datab(W_alu_result_3),
	.datac(W_alu_result_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
defparam \Equal2~2 .lut_mask = 16'h7F7F;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~1 (
	.dataa(W_alu_result_7),
	.datab(always1),
	.datac(W_alu_result_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~1_combout ),
	.cout());
defparam \always1~1 .lut_mask = 16'hEFEF;
defparam \always1~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_router_001 (
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	Equal5,
	F_pc_10,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	Equal0,
	F_pc_5,
	F_pc_3,
	Equal01,
	uav_read,
	F_pc_2,
	F_pc_4,
	F_pc_9,
	F_pc_1,
	Equal1,
	always1,
	Equal02,
	src_channel_6,
	Equal6,
	Equal2,
	Equal51,
	src_channel_5)/* synthesis synthesis_greybox=1 */;
input 	F_pc_26;
input 	F_pc_25;
input 	F_pc_24;
input 	F_pc_23;
input 	F_pc_22;
input 	F_pc_21;
input 	F_pc_20;
input 	F_pc_19;
input 	F_pc_18;
input 	F_pc_17;
input 	F_pc_16;
input 	F_pc_15;
input 	F_pc_14;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
output 	Equal5;
input 	F_pc_10;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
output 	Equal0;
input 	F_pc_5;
input 	F_pc_3;
output 	Equal01;
input 	uav_read;
input 	F_pc_2;
input 	F_pc_4;
input 	F_pc_9;
input 	F_pc_1;
output 	Equal1;
output 	always1;
output 	Equal02;
output 	src_channel_6;
output 	Equal6;
output 	Equal2;
output 	Equal51;
output 	src_channel_5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal5~0_combout ;
wire \Equal5~1_combout ;
wire \Equal5~2_combout ;
wire \Equal5~3_combout ;
wire \Equal1~0_combout ;
wire \always1~0_combout ;
wire \Equal0~2_combout ;
wire \src_channel[6]~0_combout ;
wire \src_channel[6]~1_combout ;
wire \Equal2~0_combout ;


cycloneive_lcell_comb \Equal5~4 (
	.dataa(\Equal5~0_combout ),
	.datab(\Equal5~1_combout ),
	.datac(\Equal5~2_combout ),
	.datad(\Equal5~3_combout ),
	.cin(gnd),
	.combout(Equal5),
	.cout());
defparam \Equal5~4 .lut_mask = 16'hFFFE;
defparam \Equal5~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(F_pc_10),
	.datab(F_pc_8),
	.datac(F_pc_7),
	.datad(F_pc_6),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(F_pc_5),
	.datad(F_pc_3),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h0FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(Equal5),
	.datab(Equal0),
	.datac(\Equal1~0_combout ),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hFEFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~1 (
	.dataa(Equal5),
	.datab(Equal0),
	.datac(\Equal1~0_combout ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
defparam \always1~1 .lut_mask = 16'hFFFE;
defparam \always1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\Equal0~2_combout ),
	.datab(gnd),
	.datac(F_pc_2),
	.datad(F_pc_4),
	.cin(gnd),
	.combout(Equal02),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hAFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~2 (
	.dataa(F_pc_9),
	.datab(F_pc_4),
	.datac(\Equal0~2_combout ),
	.datad(\src_channel[6]~1_combout ),
	.cin(gnd),
	.combout(src_channel_6),
	.cout());
defparam \src_channel[6]~2 .lut_mask = 16'hBFFF;
defparam \src_channel[6]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(F_pc_26),
	.datad(F_pc_25),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~0 .lut_mask = 16'h0FFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(Equal5),
	.datab(Equal0),
	.datac(Equal01),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hFFFE;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~5 (
	.dataa(Equal5),
	.datab(F_pc_10),
	.datac(gnd),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(Equal51),
	.cout());
defparam \Equal5~5 .lut_mask = 16'hEEFF;
defparam \Equal5~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[5]~3 (
	.dataa(src_channel_6),
	.datab(F_pc_26),
	.datac(F_pc_25),
	.datad(Equal02),
	.cin(gnd),
	.combout(src_channel_5),
	.cout());
defparam \src_channel[5]~3 .lut_mask = 16'hBFFF;
defparam \src_channel[5]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~0 (
	.dataa(F_pc_26),
	.datab(F_pc_25),
	.datac(F_pc_24),
	.datad(F_pc_23),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'hBFFF;
defparam \Equal5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~1 (
	.dataa(F_pc_22),
	.datab(F_pc_21),
	.datac(F_pc_20),
	.datad(F_pc_19),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
defparam \Equal5~1 .lut_mask = 16'h7FFF;
defparam \Equal5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~2 (
	.dataa(F_pc_18),
	.datab(F_pc_17),
	.datac(F_pc_16),
	.datad(F_pc_15),
	.cin(gnd),
	.combout(\Equal5~2_combout ),
	.cout());
defparam \Equal5~2 .lut_mask = 16'h7FFF;
defparam \Equal5~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~3 (
	.dataa(F_pc_14),
	.datab(F_pc_13),
	.datac(F_pc_12),
	.datad(F_pc_11),
	.cin(gnd),
	.combout(\Equal5~3_combout ),
	.cout());
defparam \Equal5~3 .lut_mask = 16'h7FFF;
defparam \Equal5~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(F_pc_2),
	.datad(F_pc_4),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hAFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(uav_read),
	.datab(F_pc_5),
	.datac(F_pc_1),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(Equal5),
	.datab(Equal0),
	.datac(Equal01),
	.datad(F_pc_9),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~0 (
	.dataa(F_pc_5),
	.datab(uav_read),
	.datac(F_pc_1),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\src_channel[6]~0_combout ),
	.cout());
defparam \src_channel[6]~0 .lut_mask = 16'hFFFD;
defparam \src_channel[6]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[6]~1 (
	.dataa(F_pc_10),
	.datab(Equal0),
	.datac(Equal5),
	.datad(\src_channel[6]~0_combout ),
	.cin(gnd),
	.combout(\src_channel[6]~1_combout ),
	.cout());
defparam \src_channel[6]~1 .lut_mask = 16'hFFFE;
defparam \src_channel[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(F_pc_4),
	.datab(F_pc_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hBBBB;
defparam \Equal2~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_router_002_5 (
	mem_86_0,
	mem_68_0,
	always0)/* synthesis synthesis_greybox=1 */;
input 	mem_86_0;
input 	mem_68_0;
output 	always0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \always0~0 (
	.dataa(mem_86_0),
	.datab(mem_68_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hEEEE;
defparam \always0~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux (
	mem_86_0,
	mem_68_0,
	in_data_toggle,
	dreg_0,
	in_data_toggle1,
	dreg_01,
	take_in_data,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	mem_86_0;
input 	mem_68_0;
input 	in_data_toggle;
input 	dreg_0;
input 	in_data_toggle1;
input 	dreg_01;
input 	take_in_data;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;


cycloneive_lcell_comb \WideOr0~1 (
	.dataa(\WideOr0~0_combout ),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(take_in_data),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hBEFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(mem_86_0),
	.datab(mem_68_0),
	.datac(in_data_toggle),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_1 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_2 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_3 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_4 (
	mem_86_0,
	mem_68_0,
	in_data_toggle,
	dreg_0,
	in_data_toggle1,
	dreg_01,
	always0,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	mem_86_0;
input 	mem_68_0;
input 	in_data_toggle;
input 	dreg_0;
input 	in_data_toggle1;
input 	dreg_01;
input 	always0;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;


cycloneive_lcell_comb \WideOr0~1 (
	.dataa(\WideOr0~0_combout ),
	.datab(in_data_toggle1),
	.datac(dreg_01),
	.datad(always0),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hBEFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(mem_86_0),
	.datab(mem_68_0),
	.datac(in_data_toggle),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEFFE;
defparam \WideOr0~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_demux_001_5 (
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_mux (
	q_a_0,
	readdata_0,
	q_a_1,
	readdata_1,
	readdata_2,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	readdata_16,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	readdata_17,
	q_a_17,
	q_a_10,
	q_a_9,
	q_a_23,
	readdata_8,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	mem_86_0,
	mem_68_0,
	src0_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid,
	out_data_toggle_flopped1,
	dreg_01,
	out_valid1,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	mem_86_01,
	mem_68_01,
	src0_valid1,
	src0_valid2,
	read_latency_shift_reg_05,
	mem_86_02,
	mem_68_02,
	src0_valid3,
	src0_valid4,
	WideOr11,
	mem_67_0,
	src_payload,
	av_readdata_pre_30,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_1,
	av_readdata_pre_11,
	av_readdata_pre_2,
	av_readdata_pre_3,
	readdata_3,
	av_readdata_pre_4,
	readdata_4,
	av_readdata_pre_111,
	av_readdata_pre_13,
	av_readdata_pre_161,
	av_readdata_pre_12,
	readdata_5,
	av_readdata_pre_5,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_211,
	av_readdata_pre_181,
	av_readdata_pre_171,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_23,
	av_readdata_pre_8,
	av_readdata_pre_221,
	readdata_7,
	av_readdata_pre_7,
	readdata_6,
	av_readdata_pre_6,
	av_readdata_pre_201,
	av_readdata_pre_191,
	src_payload1,
	av_readdata_pre_02,
	av_readdata_pre_03,
	out_data_buffer_0,
	out_data_buffer_01,
	av_readdata_pre_04,
	src_data_0,
	src_data_1,
	av_readdata_pre_110,
	av_readdata_pre_112,
	out_data_buffer_1,
	av_readdata_pre_113,
	out_data_buffer_11,
	src_data_11,
	src_data_2,
	av_readdata_pre_24,
	av_readdata_pre_25,
	out_data_buffer_2,
	av_readdata_pre_26,
	out_data_buffer_21,
	src_data_21,
	src_data_3,
	av_readdata_pre_31,
	av_readdata_pre_32,
	out_data_buffer_3,
	av_readdata_pre_33,
	out_data_buffer_31,
	src_data_31,
	src_data_4,
	av_readdata_pre_41,
	av_readdata_pre_42,
	out_data_buffer_4,
	av_readdata_pre_43,
	out_data_buffer_41,
	src_data_41,
	av_readdata_pre_51,
	av_readdata_pre_52,
	src_data_5,
	out_data_buffer_5,
	av_readdata_pre_53,
	out_data_buffer_51,
	src_data_6,
	av_readdata_pre_61,
	av_readdata_pre_62,
	out_data_buffer_6,
	av_readdata_pre_63,
	out_data_buffer_61,
	src_data_61,
	av_readdata_pre_71,
	av_readdata_pre_72,
	src_data_7,
	out_data_buffer_7,
	av_readdata_pre_73,
	out_data_buffer_71,
	out_data_buffer_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	out_data_buffer_81,
	src_data_8,
	av_readdata_pre_91,
	av_readdata_pre_92,
	out_data_buffer_9,
	out_data_buffer_91,
	src_data_9,
	out_data_buffer_10,
	av_readdata_pre_101,
	av_readdata_pre_102,
	out_data_buffer_101,
	src_data_10,
	out_data_buffer_111,
	out_data_buffer_112,
	av_readdata_pre_114,
	src_data_111,
	av_readdata_pre_121,
	av_readdata_pre_122,
	out_data_buffer_12,
	out_data_buffer_121,
	src_data_12,
	av_readdata_pre_131,
	av_readdata_pre_132,
	out_data_buffer_13,
	out_data_buffer_131,
	src_data_13,
	out_data_buffer_14,
	av_readdata_pre_141,
	av_readdata_pre_142,
	out_data_buffer_141,
	src_data_14,
	av_readdata_pre_151,
	av_readdata_pre_152,
	out_data_buffer_15,
	out_data_buffer_151,
	src_data_15,
	out_data_buffer_16,
	av_readdata_pre_162,
	out_data_buffer_161,
	src_data_16,
	out_data_buffer_17,
	out_data_buffer_171,
	av_readdata_pre_172,
	src_data_17,
	out_data_buffer_23,
	out_data_buffer_231,
	src_data_23,
	out_data_buffer_22,
	out_data_buffer_221,
	src_data_22,
	out_data_buffer_211,
	out_data_buffer_212,
	src_data_211,
	out_data_buffer_20,
	out_data_buffer_201,
	src_data_20,
	out_data_buffer_19,
	out_data_buffer_191,
	src_data_19,
	out_data_buffer_18,
	out_data_buffer_181,
	src_data_18,
	src_data_51,
	src_data_71)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	readdata_0;
input 	q_a_1;
input 	readdata_1;
input 	readdata_2;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_11;
input 	q_a_13;
input 	readdata_16;
input 	q_a_16;
input 	q_a_12;
input 	q_a_5;
input 	q_a_14;
input 	q_a_15;
input 	q_a_21;
input 	q_a_18;
input 	readdata_17;
input 	q_a_17;
input 	q_a_10;
input 	q_a_9;
input 	q_a_23;
input 	readdata_8;
input 	q_a_8;
input 	q_a_22;
input 	q_a_7;
input 	q_a_6;
input 	q_a_20;
input 	q_a_19;
input 	av_readdata_pre_16;
input 	av_readdata_pre_17;
input 	av_readdata_pre_22;
input 	av_readdata_pre_21;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_18;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	mem_86_0;
input 	mem_68_0;
input 	src0_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid;
input 	out_data_toggle_flopped1;
input 	dreg_01;
input 	out_valid1;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
input 	mem_86_01;
input 	mem_68_01;
input 	src0_valid1;
input 	src0_valid2;
input 	read_latency_shift_reg_05;
input 	mem_86_02;
input 	mem_68_02;
input 	src0_valid3;
input 	src0_valid4;
output 	WideOr11;
input 	mem_67_0;
output 	src_payload;
input 	av_readdata_pre_30;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_1;
input 	av_readdata_pre_11;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	readdata_3;
input 	av_readdata_pre_4;
input 	readdata_4;
input 	av_readdata_pre_111;
input 	av_readdata_pre_13;
input 	av_readdata_pre_161;
input 	av_readdata_pre_12;
input 	readdata_5;
input 	av_readdata_pre_5;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_211;
input 	av_readdata_pre_181;
input 	av_readdata_pre_171;
input 	av_readdata_pre_10;
input 	av_readdata_pre_9;
input 	av_readdata_pre_23;
input 	av_readdata_pre_8;
input 	av_readdata_pre_221;
input 	readdata_7;
input 	av_readdata_pre_7;
input 	readdata_6;
input 	av_readdata_pre_6;
input 	av_readdata_pre_201;
input 	av_readdata_pre_191;
output 	src_payload1;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
input 	out_data_buffer_0;
input 	out_data_buffer_01;
input 	av_readdata_pre_04;
output 	src_data_0;
output 	src_data_1;
input 	av_readdata_pre_110;
input 	av_readdata_pre_112;
input 	out_data_buffer_1;
input 	av_readdata_pre_113;
input 	out_data_buffer_11;
output 	src_data_11;
output 	src_data_2;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	out_data_buffer_2;
input 	av_readdata_pre_26;
input 	out_data_buffer_21;
output 	src_data_21;
output 	src_data_3;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
input 	out_data_buffer_3;
input 	av_readdata_pre_33;
input 	out_data_buffer_31;
output 	src_data_31;
output 	src_data_4;
input 	av_readdata_pre_41;
input 	av_readdata_pre_42;
input 	out_data_buffer_4;
input 	av_readdata_pre_43;
input 	out_data_buffer_41;
output 	src_data_41;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
output 	src_data_5;
input 	out_data_buffer_5;
input 	av_readdata_pre_53;
input 	out_data_buffer_51;
output 	src_data_6;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	out_data_buffer_6;
input 	av_readdata_pre_63;
input 	out_data_buffer_61;
output 	src_data_61;
input 	av_readdata_pre_71;
input 	av_readdata_pre_72;
output 	src_data_7;
input 	out_data_buffer_7;
input 	av_readdata_pre_73;
input 	out_data_buffer_71;
input 	out_data_buffer_8;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
input 	out_data_buffer_81;
output 	src_data_8;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
input 	out_data_buffer_9;
input 	out_data_buffer_91;
output 	src_data_9;
input 	out_data_buffer_10;
input 	av_readdata_pre_101;
input 	av_readdata_pre_102;
input 	out_data_buffer_101;
output 	src_data_10;
input 	out_data_buffer_111;
input 	out_data_buffer_112;
input 	av_readdata_pre_114;
output 	src_data_111;
input 	av_readdata_pre_121;
input 	av_readdata_pre_122;
input 	out_data_buffer_12;
input 	out_data_buffer_121;
output 	src_data_12;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
input 	out_data_buffer_13;
input 	out_data_buffer_131;
output 	src_data_13;
input 	out_data_buffer_14;
input 	av_readdata_pre_141;
input 	av_readdata_pre_142;
input 	out_data_buffer_141;
output 	src_data_14;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
input 	out_data_buffer_15;
input 	out_data_buffer_151;
output 	src_data_15;
input 	out_data_buffer_16;
input 	av_readdata_pre_162;
input 	out_data_buffer_161;
output 	src_data_16;
input 	out_data_buffer_17;
input 	out_data_buffer_171;
input 	av_readdata_pre_172;
output 	src_data_17;
input 	out_data_buffer_23;
input 	out_data_buffer_231;
output 	src_data_23;
input 	out_data_buffer_22;
input 	out_data_buffer_221;
output 	src_data_22;
input 	out_data_buffer_211;
input 	out_data_buffer_212;
output 	src_data_211;
input 	out_data_buffer_20;
input 	out_data_buffer_201;
output 	src_data_20;
input 	out_data_buffer_19;
input 	out_data_buffer_191;
output 	src_data_19;
input 	out_data_buffer_18;
input 	out_data_buffer_181;
output 	src_data_18;
output 	src_data_51;
output 	src_data_71;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;
wire \WideOr1~1_combout ;
wire \src_data[0]~4_combout ;
wire \src_data[0]~5_combout ;
wire \src_data[0]~6_combout ;
wire \src_data[0]~7_combout ;
wire \src_data[0]~8_combout ;
wire \src_data[1]~10_combout ;
wire \src_payload~2_combout ;
wire \src_data[1]~12_combout ;
wire \src_data[1]~13_combout ;
wire \src_data[2]~15_combout ;
wire \src_data[2]~17_combout ;
wire \src_data[2]~18_combout ;
wire \src_data[3]~20_combout ;
wire \src_data[3]~22_combout ;
wire \src_data[3]~23_combout ;
wire \src_data[4]~25_combout ;
wire \src_data[4]~27_combout ;
wire \src_data[4]~28_combout ;
wire \src_data[5]~30_combout ;
wire \src_data[5]~31_combout ;
wire \src_data[6]~34_combout ;
wire \src_data[6]~36_combout ;
wire \src_data[6]~37_combout ;
wire \src_data[7]~39_combout ;
wire \src_data[7]~40_combout ;
wire \src_payload~3_combout ;
wire \src_data[8]~43_combout ;
wire \src_data[8]~44_combout ;
wire \src_data[8]~45_combout ;
wire \src_data[9]~46_combout ;
wire \src_data[9]~47_combout ;
wire \src_data[9]~48_combout ;
wire \src_data[10]~49_combout ;
wire \src_data[10]~50_combout ;
wire \src_data[10]~51_combout ;
wire \src_data[11]~52_combout ;
wire \src_data[11]~53_combout ;
wire \src_data[12]~54_combout ;
wire \src_data[12]~55_combout ;
wire \src_data[12]~56_combout ;
wire \src_data[13]~57_combout ;
wire \src_data[13]~58_combout ;
wire \src_data[13]~59_combout ;
wire \src_data[14]~60_combout ;
wire \src_data[14]~61_combout ;
wire \src_data[14]~62_combout ;
wire \src_data[15]~63_combout ;
wire \src_data[15]~64_combout ;
wire \src_data[15]~65_combout ;
wire \src_payload~4_combout ;
wire \src_data[16]~66_combout ;
wire \src_data[16]~67_combout ;
wire \src_data[16]~68_combout ;
wire \src_data[17]~69_combout ;
wire \src_data[17]~70_combout ;
wire \src_payload~5_combout ;
wire \src_data[17]~71_combout ;
wire \src_data[23]~72_combout ;
wire \src_payload~6_combout ;
wire \src_data[22]~74_combout ;
wire \src_data[22]~75_combout ;
wire \src_payload~7_combout ;
wire \src_data[21]~76_combout ;
wire \src_data[21]~77_combout ;
wire \src_data[20]~78_combout ;
wire \src_data[20]~79_combout ;
wire \src_data[19]~80_combout ;
wire \src_data[19]~81_combout ;
wire \src_data[18]~82_combout ;
wire \src_data[18]~83_combout ;
wire \src_payload~8_combout ;
wire \src_data[5]~33_combout ;
wire \src_data[7]~42_combout ;


cycloneive_lcell_comb WideOr1(
	.dataa(\WideOr1~0_combout ),
	.datab(\WideOr1~1_combout ),
	.datac(src0_valid3),
	.datad(src0_valid4),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_02),
	.datab(mem_67_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_04),
	.datab(av_readdata_pre_30),
	.datac(mem_86_01),
	.datad(mem_68_01),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEFFF;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~9 (
	.dataa(\src_data[0]~5_combout ),
	.datab(\src_data[0]~8_combout ),
	.datac(read_latency_shift_reg_02),
	.datad(av_readdata_pre_04),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0]~9 .lut_mask = 16'hFFFE;
defparam \src_data[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~11 (
	.dataa(\src_data[1]~10_combout ),
	.datab(\src_payload~2_combout ),
	.datac(src0_valid4),
	.datad(q_a_1),
	.cin(gnd),
	.combout(src_data_1),
	.cout());
defparam \src_data[1]~11 .lut_mask = 16'hFFFE;
defparam \src_data[1]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~14 (
	.dataa(\src_data[1]~12_combout ),
	.datab(\src_data[1]~13_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_11),
	.cin(gnd),
	.combout(src_data_11),
	.cout());
defparam \src_data[1]~14 .lut_mask = 16'hFFFE;
defparam \src_data[1]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~16 (
	.dataa(src_payload1),
	.datab(\src_data[2]~15_combout ),
	.datac(src0_valid),
	.datad(readdata_2),
	.cin(gnd),
	.combout(src_data_2),
	.cout());
defparam \src_data[2]~16 .lut_mask = 16'hFFFE;
defparam \src_data[2]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~19 (
	.dataa(\src_data[2]~17_combout ),
	.datab(\src_data[2]~18_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_21),
	.cin(gnd),
	.combout(src_data_21),
	.cout());
defparam \src_data[2]~19 .lut_mask = 16'hFFFE;
defparam \src_data[2]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~21 (
	.dataa(src_payload1),
	.datab(\src_data[3]~20_combout ),
	.datac(src0_valid),
	.datad(readdata_3),
	.cin(gnd),
	.combout(src_data_3),
	.cout());
defparam \src_data[3]~21 .lut_mask = 16'hFFFE;
defparam \src_data[3]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~24 (
	.dataa(\src_data[3]~22_combout ),
	.datab(\src_data[3]~23_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_31),
	.cin(gnd),
	.combout(src_data_31),
	.cout());
defparam \src_data[3]~24 .lut_mask = 16'hFFFE;
defparam \src_data[3]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~26 (
	.dataa(src_payload1),
	.datab(\src_data[4]~25_combout ),
	.datac(src0_valid),
	.datad(readdata_4),
	.cin(gnd),
	.combout(src_data_4),
	.cout());
defparam \src_data[4]~26 .lut_mask = 16'hFFFE;
defparam \src_data[4]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~29 (
	.dataa(\src_data[4]~27_combout ),
	.datab(\src_data[4]~28_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_41),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[4]~29 .lut_mask = 16'hFFFE;
defparam \src_data[4]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~32 (
	.dataa(\src_data[5]~30_combout ),
	.datab(\src_data[5]~31_combout ),
	.datac(src0_valid4),
	.datad(q_a_5),
	.cin(gnd),
	.combout(src_data_5),
	.cout());
defparam \src_data[5]~32 .lut_mask = 16'hFFFE;
defparam \src_data[5]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~35 (
	.dataa(src_payload1),
	.datab(\src_data[6]~34_combout ),
	.datac(src0_valid),
	.datad(readdata_6),
	.cin(gnd),
	.combout(src_data_6),
	.cout());
defparam \src_data[6]~35 .lut_mask = 16'hFFFE;
defparam \src_data[6]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~38 (
	.dataa(\src_data[6]~36_combout ),
	.datab(\src_data[6]~37_combout ),
	.datac(out_valid),
	.datad(out_data_buffer_61),
	.cin(gnd),
	.combout(src_data_61),
	.cout());
defparam \src_data[6]~38 .lut_mask = 16'hFFFE;
defparam \src_data[6]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~41 (
	.dataa(\src_data[7]~39_combout ),
	.datab(\src_data[7]~40_combout ),
	.datac(src0_valid4),
	.datad(q_a_7),
	.cin(gnd),
	.combout(src_data_7),
	.cout());
defparam \src_data[7]~41 .lut_mask = 16'hFFFE;
defparam \src_data[7]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8] (
	.dataa(\src_data[8]~44_combout ),
	.datab(\src_data[8]~45_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_81),
	.cin(gnd),
	.combout(src_data_8),
	.cout());
defparam \src_data[8] .lut_mask = 16'hFFFE;
defparam \src_data[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9] (
	.dataa(\src_data[9]~46_combout ),
	.datab(\src_data[9]~47_combout ),
	.datac(\src_data[9]~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_9),
	.cout());
defparam \src_data[9] .lut_mask = 16'hFEFE;
defparam \src_data[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10] (
	.dataa(\src_data[10]~50_combout ),
	.datab(\src_data[10]~51_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_101),
	.cin(gnd),
	.combout(src_data_10),
	.cout());
defparam \src_data[10] .lut_mask = 16'hFFFE;
defparam \src_data[10] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11] (
	.dataa(\src_data[11]~52_combout ),
	.datab(\src_data[11]~53_combout ),
	.datac(read_latency_shift_reg_03),
	.datad(av_readdata_pre_114),
	.cin(gnd),
	.combout(src_data_111),
	.cout());
defparam \src_data[11] .lut_mask = 16'hFFFE;
defparam \src_data[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12] (
	.dataa(\src_data[12]~54_combout ),
	.datab(\src_data[12]~55_combout ),
	.datac(\src_data[12]~56_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_12),
	.cout());
defparam \src_data[12] .lut_mask = 16'hFEFE;
defparam \src_data[12] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13] (
	.dataa(\src_data[13]~57_combout ),
	.datab(\src_data[13]~58_combout ),
	.datac(\src_data[13]~59_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_13),
	.cout());
defparam \src_data[13] .lut_mask = 16'hFEFE;
defparam \src_data[13] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14] (
	.dataa(\src_data[14]~61_combout ),
	.datab(\src_data[14]~62_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_141),
	.cin(gnd),
	.combout(src_data_14),
	.cout());
defparam \src_data[14] .lut_mask = 16'hFFFE;
defparam \src_data[14] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15] (
	.dataa(\src_data[15]~63_combout ),
	.datab(\src_data[15]~64_combout ),
	.datac(\src_data[15]~65_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_15),
	.cout());
defparam \src_data[15] .lut_mask = 16'hFEFE;
defparam \src_data[15] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16] (
	.dataa(\src_data[16]~67_combout ),
	.datab(\src_data[16]~68_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_161),
	.cin(gnd),
	.combout(src_data_16),
	.cout());
defparam \src_data[16] .lut_mask = 16'hFFFE;
defparam \src_data[16] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17] (
	.dataa(\src_data[17]~69_combout ),
	.datab(\src_data[17]~70_combout ),
	.datac(\src_payload~5_combout ),
	.datad(\src_data[17]~71_combout ),
	.cin(gnd),
	.combout(src_data_17),
	.cout());
defparam \src_data[17] .lut_mask = 16'hFFFE;
defparam \src_data[17] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~73 (
	.dataa(\src_data[23]~72_combout ),
	.datab(\src_payload~6_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_231),
	.cin(gnd),
	.combout(src_data_23),
	.cout());
defparam \src_data[23]~73 .lut_mask = 16'hFFFE;
defparam \src_data[23]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22] (
	.dataa(\src_data[22]~75_combout ),
	.datab(\src_payload~7_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_221),
	.cin(gnd),
	.combout(src_data_22),
	.cout());
defparam \src_data[22] .lut_mask = 16'hFFFE;
defparam \src_data[22] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21] (
	.dataa(\src_data[21]~76_combout ),
	.datab(\src_data[21]~77_combout ),
	.datac(read_latency_shift_reg_0),
	.datad(av_readdata_pre_21),
	.cin(gnd),
	.combout(src_data_211),
	.cout());
defparam \src_data[21] .lut_mask = 16'hFFFE;
defparam \src_data[21] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20] (
	.dataa(\src_data[20]~78_combout ),
	.datab(\src_data[20]~79_combout ),
	.datac(read_latency_shift_reg_0),
	.datad(av_readdata_pre_20),
	.cin(gnd),
	.combout(src_data_20),
	.cout());
defparam \src_data[20] .lut_mask = 16'hFFFE;
defparam \src_data[20] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19] (
	.dataa(\src_data[19]~80_combout ),
	.datab(\src_data[19]~81_combout ),
	.datac(read_latency_shift_reg_0),
	.datad(av_readdata_pre_19),
	.cin(gnd),
	.combout(src_data_19),
	.cout());
defparam \src_data[19] .lut_mask = 16'hFFFE;
defparam \src_data[19] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18] (
	.dataa(\src_data[18]~83_combout ),
	.datab(\src_payload~8_combout ),
	.datac(out_valid1),
	.datad(out_data_buffer_181),
	.cin(gnd),
	.combout(src_data_18),
	.cout());
defparam \src_data[18] .lut_mask = 16'hFFFE;
defparam \src_data[18] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~84 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[5]~33_combout ),
	.datad(out_data_buffer_51),
	.cin(gnd),
	.combout(src_data_51),
	.cout());
defparam \src_data[5]~84 .lut_mask = 16'hFFF6;
defparam \src_data[5]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~85 (
	.dataa(out_data_toggle_flopped),
	.datab(dreg_0),
	.datac(\src_data[7]~42_combout ),
	.datad(out_data_buffer_71),
	.cin(gnd),
	.combout(src_data_71),
	.cout());
defparam \src_data[7]~85 .lut_mask = 16'hFFF6;
defparam \src_data[7]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(src0_valid),
	.datac(out_valid),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~1 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(src0_valid1),
	.datad(src0_valid2),
	.cin(gnd),
	.combout(\WideOr1~1_combout ),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'hFFFE;
defparam \WideOr1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~4 (
	.dataa(src0_valid2),
	.datab(src0_valid3),
	.datac(av_readdata_pre_01),
	.datad(av_readdata_pre_0),
	.cin(gnd),
	.combout(\src_data[0]~4_combout ),
	.cout());
defparam \src_data[0]~4 .lut_mask = 16'hFFFE;
defparam \src_data[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~5 (
	.dataa(src_payload1),
	.datab(\src_data[0]~4_combout ),
	.datac(src0_valid),
	.datad(readdata_0),
	.cin(gnd),
	.combout(\src_data[0]~5_combout ),
	.cout());
defparam \src_data[0]~5 .lut_mask = 16'hFFFE;
defparam \src_data[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~6 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_02),
	.datad(av_readdata_pre_03),
	.cin(gnd),
	.combout(\src_data[0]~6_combout ),
	.cout());
defparam \src_data[0]~6 .lut_mask = 16'hFFFE;
defparam \src_data[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~7 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_0),
	.datad(out_data_buffer_01),
	.cin(gnd),
	.combout(\src_data[0]~7_combout ),
	.cout());
defparam \src_data[0]~7 .lut_mask = 16'hFFFE;
defparam \src_data[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~8 (
	.dataa(\src_data[0]~6_combout ),
	.datab(\src_data[0]~7_combout ),
	.datac(src0_valid4),
	.datad(q_a_0),
	.cin(gnd),
	.combout(\src_data[0]~8_combout ),
	.cout());
defparam \src_data[0]~8 .lut_mask = 16'hFFFE;
defparam \src_data[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~10 (
	.dataa(src0_valid),
	.datab(src0_valid2),
	.datac(av_readdata_pre_1),
	.datad(readdata_1),
	.cin(gnd),
	.combout(\src_data[1]~10_combout ),
	.cout());
defparam \src_data[1]~10 .lut_mask = 16'hFFFE;
defparam \src_data[1]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_05),
	.datab(av_readdata_pre_11),
	.datac(mem_86_02),
	.datad(mem_68_02),
	.cin(gnd),
	.combout(\src_payload~2_combout ),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEFFF;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~12 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_110),
	.datad(av_readdata_pre_112),
	.cin(gnd),
	.combout(\src_data[1]~12_combout ),
	.cout());
defparam \src_data[1]~12 .lut_mask = 16'hFFFE;
defparam \src_data[1]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~13 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_1),
	.datad(av_readdata_pre_113),
	.cin(gnd),
	.combout(\src_data[1]~13_combout ),
	.cout());
defparam \src_data[1]~13 .lut_mask = 16'hFFFE;
defparam \src_data[1]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~15 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_2),
	.datad(av_readdata_pre_2),
	.cin(gnd),
	.combout(\src_data[2]~15_combout ),
	.cout());
defparam \src_data[2]~15 .lut_mask = 16'hFFFE;
defparam \src_data[2]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~17 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_24),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\src_data[2]~17_combout ),
	.cout());
defparam \src_data[2]~17 .lut_mask = 16'hFFFE;
defparam \src_data[2]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~18 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_2),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\src_data[2]~18_combout ),
	.cout());
defparam \src_data[2]~18 .lut_mask = 16'hFFFE;
defparam \src_data[2]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~20 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_3),
	.datad(av_readdata_pre_3),
	.cin(gnd),
	.combout(\src_data[3]~20_combout ),
	.cout());
defparam \src_data[3]~20 .lut_mask = 16'hFFFE;
defparam \src_data[3]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~22 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_31),
	.datad(av_readdata_pre_32),
	.cin(gnd),
	.combout(\src_data[3]~22_combout ),
	.cout());
defparam \src_data[3]~22 .lut_mask = 16'hFFFE;
defparam \src_data[3]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~23 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_3),
	.datad(av_readdata_pre_33),
	.cin(gnd),
	.combout(\src_data[3]~23_combout ),
	.cout());
defparam \src_data[3]~23 .lut_mask = 16'hFFFE;
defparam \src_data[3]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~25 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_4),
	.datad(av_readdata_pre_4),
	.cin(gnd),
	.combout(\src_data[4]~25_combout ),
	.cout());
defparam \src_data[4]~25 .lut_mask = 16'hFFFE;
defparam \src_data[4]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~27 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_41),
	.datad(av_readdata_pre_42),
	.cin(gnd),
	.combout(\src_data[4]~27_combout ),
	.cout());
defparam \src_data[4]~27 .lut_mask = 16'hFFFE;
defparam \src_data[4]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~28 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_4),
	.datad(av_readdata_pre_43),
	.cin(gnd),
	.combout(\src_data[4]~28_combout ),
	.cout());
defparam \src_data[4]~28 .lut_mask = 16'hFFFE;
defparam \src_data[4]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~30 (
	.dataa(src0_valid),
	.datab(src0_valid2),
	.datac(av_readdata_pre_5),
	.datad(readdata_5),
	.cin(gnd),
	.combout(\src_data[5]~30_combout ),
	.cout());
defparam \src_data[5]~30 .lut_mask = 16'hFFFE;
defparam \src_data[5]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~31 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_51),
	.datad(av_readdata_pre_52),
	.cin(gnd),
	.combout(\src_data[5]~31_combout ),
	.cout());
defparam \src_data[5]~31 .lut_mask = 16'hFFFE;
defparam \src_data[5]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~34 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_6),
	.datad(av_readdata_pre_6),
	.cin(gnd),
	.combout(\src_data[6]~34_combout ),
	.cout());
defparam \src_data[6]~34 .lut_mask = 16'hFFFE;
defparam \src_data[6]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~36 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_61),
	.datad(av_readdata_pre_62),
	.cin(gnd),
	.combout(\src_data[6]~36_combout ),
	.cout());
defparam \src_data[6]~36 .lut_mask = 16'hFFFE;
defparam \src_data[6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~37 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_6),
	.datad(av_readdata_pre_63),
	.cin(gnd),
	.combout(\src_data[6]~37_combout ),
	.cout());
defparam \src_data[6]~37 .lut_mask = 16'hFFFE;
defparam \src_data[6]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~39 (
	.dataa(src0_valid),
	.datab(src0_valid2),
	.datac(av_readdata_pre_7),
	.datad(readdata_7),
	.cin(gnd),
	.combout(\src_data[7]~39_combout ),
	.cout());
defparam \src_data[7]~39 .lut_mask = 16'hFFFE;
defparam \src_data[7]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~40 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_71),
	.datad(av_readdata_pre_72),
	.cin(gnd),
	.combout(\src_data[7]~40_combout ),
	.cout());
defparam \src_data[7]~40 .lut_mask = 16'hFFFE;
defparam \src_data[7]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_01),
	.datab(readdata_8),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(\src_payload~3_combout ),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEFFF;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~43 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_8),
	.datad(out_data_buffer_8),
	.cin(gnd),
	.combout(\src_data[8]~43_combout ),
	.cout());
defparam \src_data[8]~43 .lut_mask = 16'hFFFE;
defparam \src_data[8]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~44 (
	.dataa(\src_payload~3_combout ),
	.datab(\src_data[8]~43_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_8),
	.cin(gnd),
	.combout(\src_data[8]~44_combout ),
	.cout());
defparam \src_data[8]~44 .lut_mask = 16'hFFFE;
defparam \src_data[8]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~45 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_81),
	.datad(av_readdata_pre_82),
	.cin(gnd),
	.combout(\src_data[8]~45_combout ),
	.cout());
defparam \src_data[8]~45 .lut_mask = 16'hFFFE;
defparam \src_data[8]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~46 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_91),
	.datad(av_readdata_pre_92),
	.cin(gnd),
	.combout(\src_data[9]~46_combout ),
	.cout());
defparam \src_data[9]~46 .lut_mask = 16'hFFFE;
defparam \src_data[9]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~47 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_9),
	.datad(av_readdata_pre_9),
	.cin(gnd),
	.combout(\src_data[9]~47_combout ),
	.cout());
defparam \src_data[9]~47 .lut_mask = 16'hFFFE;
defparam \src_data[9]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~48 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_9),
	.datad(out_data_buffer_91),
	.cin(gnd),
	.combout(\src_data[9]~48_combout ),
	.cout());
defparam \src_data[9]~48 .lut_mask = 16'hFFFE;
defparam \src_data[9]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~49 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_10),
	.datad(out_data_buffer_10),
	.cin(gnd),
	.combout(\src_data[10]~49_combout ),
	.cout());
defparam \src_data[10]~49 .lut_mask = 16'hFFFE;
defparam \src_data[10]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~50 (
	.dataa(src_payload1),
	.datab(\src_data[10]~49_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\src_data[10]~50_combout ),
	.cout());
defparam \src_data[10]~50 .lut_mask = 16'hFFFE;
defparam \src_data[10]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~51 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_101),
	.datad(av_readdata_pre_102),
	.cin(gnd),
	.combout(\src_data[10]~51_combout ),
	.cout());
defparam \src_data[10]~51 .lut_mask = 16'hFFFE;
defparam \src_data[10]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~52 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_11),
	.datad(av_readdata_pre_111),
	.cin(gnd),
	.combout(\src_data[11]~52_combout ),
	.cout());
defparam \src_data[11]~52 .lut_mask = 16'hFFFE;
defparam \src_data[11]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~53 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_111),
	.datad(out_data_buffer_112),
	.cin(gnd),
	.combout(\src_data[11]~53_combout ),
	.cout());
defparam \src_data[11]~53 .lut_mask = 16'hFFFE;
defparam \src_data[11]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~54 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_121),
	.datad(av_readdata_pre_122),
	.cin(gnd),
	.combout(\src_data[12]~54_combout ),
	.cout());
defparam \src_data[12]~54 .lut_mask = 16'hFFFE;
defparam \src_data[12]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~55 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_12),
	.datad(av_readdata_pre_12),
	.cin(gnd),
	.combout(\src_data[12]~55_combout ),
	.cout());
defparam \src_data[12]~55 .lut_mask = 16'hFFFE;
defparam \src_data[12]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~56 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_12),
	.datad(out_data_buffer_121),
	.cin(gnd),
	.combout(\src_data[12]~56_combout ),
	.cout());
defparam \src_data[12]~56 .lut_mask = 16'hFFFE;
defparam \src_data[12]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~57 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_131),
	.datad(av_readdata_pre_132),
	.cin(gnd),
	.combout(\src_data[13]~57_combout ),
	.cout());
defparam \src_data[13]~57 .lut_mask = 16'hFFFE;
defparam \src_data[13]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~58 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_13),
	.datad(av_readdata_pre_13),
	.cin(gnd),
	.combout(\src_data[13]~58_combout ),
	.cout());
defparam \src_data[13]~58 .lut_mask = 16'hFFFE;
defparam \src_data[13]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~59 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_13),
	.datad(out_data_buffer_131),
	.cin(gnd),
	.combout(\src_data[13]~59_combout ),
	.cout());
defparam \src_data[13]~59 .lut_mask = 16'hFFFE;
defparam \src_data[13]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~60 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_14),
	.datad(out_data_buffer_14),
	.cin(gnd),
	.combout(\src_data[14]~60_combout ),
	.cout());
defparam \src_data[14]~60 .lut_mask = 16'hFFFE;
defparam \src_data[14]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~61 (
	.dataa(src_payload1),
	.datab(\src_data[14]~60_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\src_data[14]~61_combout ),
	.cout());
defparam \src_data[14]~61 .lut_mask = 16'hFFFE;
defparam \src_data[14]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~62 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_141),
	.datad(av_readdata_pre_142),
	.cin(gnd),
	.combout(\src_data[14]~62_combout ),
	.cout());
defparam \src_data[14]~62 .lut_mask = 16'hFFFE;
defparam \src_data[14]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~63 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_151),
	.datad(av_readdata_pre_152),
	.cin(gnd),
	.combout(\src_data[15]~63_combout ),
	.cout());
defparam \src_data[15]~63 .lut_mask = 16'hFFFE;
defparam \src_data[15]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~64 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_15),
	.datad(av_readdata_pre_15),
	.cin(gnd),
	.combout(\src_data[15]~64_combout ),
	.cout());
defparam \src_data[15]~64 .lut_mask = 16'hFFFE;
defparam \src_data[15]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~65 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_15),
	.datad(out_data_buffer_151),
	.cin(gnd),
	.combout(\src_data[15]~65_combout ),
	.cout());
defparam \src_data[15]~65 .lut_mask = 16'hFFFE;
defparam \src_data[15]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_01),
	.datab(readdata_16),
	.datac(mem_86_0),
	.datad(mem_68_0),
	.cin(gnd),
	.combout(\src_payload~4_combout ),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEFFF;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~66 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_16),
	.datad(out_data_buffer_16),
	.cin(gnd),
	.combout(\src_data[16]~66_combout ),
	.cout());
defparam \src_data[16]~66 .lut_mask = 16'hFFFE;
defparam \src_data[16]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~67 (
	.dataa(\src_payload~4_combout ),
	.datab(\src_data[16]~66_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_161),
	.cin(gnd),
	.combout(\src_data[16]~67_combout ),
	.cout());
defparam \src_data[16]~67 .lut_mask = 16'hFFFE;
defparam \src_data[16]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~68 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_162),
	.datad(av_readdata_pre_16),
	.cin(gnd),
	.combout(\src_data[16]~68_combout ),
	.cout());
defparam \src_data[16]~68 .lut_mask = 16'hFFFE;
defparam \src_data[16]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~69 (
	.dataa(src0_valid),
	.datab(src0_valid2),
	.datac(av_readdata_pre_171),
	.datad(readdata_17),
	.cin(gnd),
	.combout(\src_data[17]~69_combout ),
	.cout());
defparam \src_data[17]~69 .lut_mask = 16'hFFFE;
defparam \src_data[17]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~70 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_17),
	.datad(out_data_buffer_17),
	.cin(gnd),
	.combout(\src_data[17]~70_combout ),
	.cout());
defparam \src_data[17]~70 .lut_mask = 16'hFFFE;
defparam \src_data[17]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(out_data_buffer_171),
	.datab(gnd),
	.datac(out_data_toggle_flopped1),
	.datad(dreg_01),
	.cin(gnd),
	.combout(\src_payload~5_combout ),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hAFFA;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~71 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_172),
	.datad(av_readdata_pre_17),
	.cin(gnd),
	.combout(\src_data[17]~71_combout ),
	.cout());
defparam \src_data[17]~71 .lut_mask = 16'hFFFE;
defparam \src_data[17]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~72 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_23),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\src_data[23]~72_combout ),
	.cout());
defparam \src_data[23]~72 .lut_mask = 16'hFFFE;
defparam \src_data[23]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(out_data_buffer_23),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\src_payload~6_combout ),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hAFFA;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~74 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_22),
	.datad(out_data_buffer_22),
	.cin(gnd),
	.combout(\src_data[22]~74_combout ),
	.cout());
defparam \src_data[22]~74 .lut_mask = 16'hFFFE;
defparam \src_data[22]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~75 (
	.dataa(src_payload1),
	.datab(\src_data[22]~74_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_221),
	.cin(gnd),
	.combout(\src_data[22]~75_combout ),
	.cout());
defparam \src_data[22]~75 .lut_mask = 16'hFFFE;
defparam \src_data[22]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~7_combout ),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~76 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_21),
	.datad(av_readdata_pre_211),
	.cin(gnd),
	.combout(\src_data[21]~76_combout ),
	.cout());
defparam \src_data[21]~76 .lut_mask = 16'hFFFE;
defparam \src_data[21]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~77 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_211),
	.datad(out_data_buffer_212),
	.cin(gnd),
	.combout(\src_data[21]~77_combout ),
	.cout());
defparam \src_data[21]~77 .lut_mask = 16'hFFFE;
defparam \src_data[21]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~78 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_20),
	.datad(av_readdata_pre_201),
	.cin(gnd),
	.combout(\src_data[20]~78_combout ),
	.cout());
defparam \src_data[20]~78 .lut_mask = 16'hFFFE;
defparam \src_data[20]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~79 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_20),
	.datad(out_data_buffer_201),
	.cin(gnd),
	.combout(\src_data[20]~79_combout ),
	.cout());
defparam \src_data[20]~79 .lut_mask = 16'hFFFE;
defparam \src_data[20]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~80 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_19),
	.datad(av_readdata_pre_191),
	.cin(gnd),
	.combout(\src_data[19]~80_combout ),
	.cout());
defparam \src_data[19]~80 .lut_mask = 16'hFFFE;
defparam \src_data[19]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~81 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_19),
	.datad(out_data_buffer_191),
	.cin(gnd),
	.combout(\src_data[19]~81_combout ),
	.cout());
defparam \src_data[19]~81 .lut_mask = 16'hFFFE;
defparam \src_data[19]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~82 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_18),
	.datad(out_data_buffer_18),
	.cin(gnd),
	.combout(\src_data[18]~82_combout ),
	.cout());
defparam \src_data[18]~82 .lut_mask = 16'hFFFE;
defparam \src_data[18]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~83 (
	.dataa(src_payload1),
	.datab(\src_data[18]~82_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_181),
	.cin(gnd),
	.combout(\src_data[18]~83_combout ),
	.cout());
defparam \src_data[18]~83 .lut_mask = 16'hFFFE;
defparam \src_data[18]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(read_latency_shift_reg_0),
	.datab(av_readdata_pre_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~8_combout ),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~33 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_5),
	.datad(av_readdata_pre_53),
	.cin(gnd),
	.combout(\src_data[5]~33_combout ),
	.cout());
defparam \src_data[5]~33 .lut_mask = 16'hFFFE;
defparam \src_data[5]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~42 (
	.dataa(read_latency_shift_reg_02),
	.datab(out_valid1),
	.datac(out_data_buffer_7),
	.datad(av_readdata_pre_73),
	.cin(gnd),
	.combout(\src_data[7]~42_combout ),
	.cout());
defparam \src_data[7]~42 .lut_mask = 16'hFFFE;
defparam \src_data[7]~42 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_mm_interconnect_0_rsp_mux_001 (
	readdata_16,
	read_latency_shift_reg_0,
	mem_86_0,
	mem_68_0,
	read_latency_shift_reg_01,
	mem_86_01,
	mem_68_01,
	read_latency_shift_reg_02,
	mem_86_02,
	mem_68_02,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src_payload,
	src_payload1,
	out_valid,
	out_valid1,
	WideOr11,
	av_readdata_pre_30,
	src_payload2,
	src_payload3,
	readdata_5,
	src_payload4)/* synthesis synthesis_greybox=1 */;
input 	readdata_16;
input 	read_latency_shift_reg_0;
input 	mem_86_0;
input 	mem_68_0;
input 	read_latency_shift_reg_01;
input 	mem_86_01;
input 	mem_68_01;
input 	read_latency_shift_reg_02;
input 	mem_86_02;
input 	mem_68_02;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
output 	src_payload;
output 	src_payload1;
input 	out_valid;
input 	out_valid1;
output 	WideOr11;
input 	av_readdata_pre_30;
output 	src_payload2;
output 	src_payload3;
input 	readdata_5;
output 	src_payload4;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;


cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_02),
	.datab(mem_86_02),
	.datac(mem_68_02),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hFEFE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_86_01),
	.datac(mem_68_01),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hFEFE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(\WideOr1~0_combout ),
	.datab(src_payload1),
	.datac(out_valid),
	.datad(out_valid1),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_86_01),
	.datac(mem_68_01),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hFFFE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(readdata_16),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hFFFE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(readdata_5),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hFFFE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(src1_valid2),
	.datad(src_payload),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0 (
	sr_0,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_11,
	W_alu_result_2,
	W_alu_result_3,
	q_a_0,
	readdata_0,
	q_a_1,
	readdata_1,
	readdata_2,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	readdata_17,
	q_a_17,
	q_a_31,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_10,
	q_a_24,
	q_a_9,
	q_a_23,
	readdata_8,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	readdata_01,
	readdata_11,
	readdata_21,
	readdata_3,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	ir_out_0,
	ir_out_1,
	d_read,
	d_write,
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_3,
	i_read,
	F_pc_2,
	F_pc_4,
	F_pc_9,
	d_writedata_0,
	d_byteenable_0,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	mem_86_0,
	mem_68_0,
	src0_valid,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	src0_valid1,
	src0_valid2,
	read_latency_shift_reg_04,
	mem_86_01,
	mem_68_01,
	src0_valid3,
	src0_valid4,
	WideOr1,
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	mem_67_04,
	mem_67_05,
	mem_67_06,
	out_data_buffer_67,
	out_data_buffer_671,
	mem_67_07,
	src_payload,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src_payload1,
	src_payload2,
	out_valid2,
	out_valid3,
	av_readdatavalid,
	WideOr11,
	local_read,
	hbreak_enabled,
	av_readdata_pre_30,
	src_payload3,
	av_readdata_pre_0,
	av_readdata_pre_01,
	out_data_buffer_0,
	out_data_buffer_01,
	av_readdata_pre_1,
	out_data_buffer_1,
	av_readdata_pre_11,
	out_data_buffer_11,
	av_readdata_pre_2,
	out_data_buffer_2,
	out_data_buffer_21,
	av_readdata_pre_3,
	readdata_31,
	out_data_buffer_3,
	out_data_buffer_31,
	av_readdata_pre_4,
	readdata_4,
	out_data_buffer_4,
	out_data_buffer_41,
	d_byteenable_2,
	mem,
	src_data_46,
	av_readdata_pre_111,
	out_data_buffer_111,
	out_data_buffer_112,
	av_readdata_pre_13,
	out_data_buffer_13,
	out_data_buffer_131,
	src_payload4,
	av_readdata_pre_16,
	out_data_buffer_16,
	out_data_buffer_161,
	av_readdata_pre_12,
	out_data_buffer_12,
	out_data_buffer_121,
	src_payload5,
	av_readdata_pre_5,
	out_data_buffer_5,
	out_data_buffer_51,
	out_data_buffer_14,
	av_readdata_pre_14,
	out_data_buffer_141,
	av_readdata_pre_15,
	out_data_buffer_15,
	out_data_buffer_151,
	av_readdata_pre_21,
	out_data_buffer_211,
	out_data_buffer_212,
	out_data_buffer_18,
	av_readdata_pre_18,
	out_data_buffer_181,
	av_readdata_pre_17,
	out_data_buffer_17,
	out_data_buffer_171,
	av_readdata_pre_31,
	out_data_buffer_311,
	out_data_buffer_312,
	out_data_buffer_30,
	av_readdata_pre_301,
	out_data_buffer_301,
	av_readdata_pre_29,
	out_data_buffer_29,
	out_data_buffer_291,
	out_data_buffer_28,
	av_readdata_pre_28,
	out_data_buffer_281,
	av_readdata_pre_27,
	out_data_buffer_27,
	out_data_buffer_271,
	out_data_buffer_26,
	av_readdata_pre_26,
	out_data_buffer_261,
	av_readdata_pre_25,
	out_data_buffer_25,
	out_data_buffer_251,
	out_data_buffer_10,
	av_readdata_pre_10,
	out_data_buffer_101,
	out_data_buffer_24,
	av_readdata_pre_24,
	out_data_buffer_241,
	av_readdata_pre_9,
	out_data_buffer_9,
	out_data_buffer_91,
	av_readdata_pre_23,
	out_data_buffer_23,
	out_data_buffer_231,
	out_data_buffer_8,
	av_readdata_pre_8,
	out_data_buffer_81,
	out_data_buffer_22,
	av_readdata_pre_22,
	out_data_buffer_221,
	readdata_7,
	out_data_buffer_7,
	av_readdata_pre_7,
	out_data_buffer_71,
	readdata_6,
	av_readdata_pre_6,
	out_data_buffer_6,
	out_data_buffer_61,
	av_readdata_pre_20,
	out_data_buffer_20,
	out_data_buffer_201,
	av_readdata_pre_19,
	out_data_buffer_19,
	out_data_buffer_191,
	src_payload6,
	src_data_0,
	av_readdata_9,
	av_readdata_8,
	dreg_1,
	r_early_rst,
	readdata_41,
	src_data_1,
	src_data_11,
	src_data_2,
	src_data_21,
	src_data_3,
	src_data_31,
	src_data_4,
	src_data_41,
	src_data_5,
	src_data_6,
	src_data_61,
	src_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_111,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	d_byteenable_1,
	d_byteenable_3,
	readdata_111,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	out_data_buffer_282,
	out_data_buffer_283,
	readdata_211,
	d_writedata_21,
	d_writedata_18,
	readdata_18,
	out_data_buffer_272,
	out_data_buffer_273,
	readdata_171,
	readdata_311,
	out_data_buffer_262,
	out_data_buffer_263,
	readdata_30,
	out_data_buffer_252,
	out_data_buffer_253,
	readdata_29,
	out_data_buffer_242,
	out_data_buffer_243,
	readdata_28,
	src_data_23,
	readdata_27,
	src_data_22,
	readdata_26,
	src_data_211,
	readdata_25,
	src_data_20,
	readdata_10,
	readdata_24,
	src_data_19,
	readdata_9,
	d_writedata_23,
	readdata_23,
	src_data_18,
	readdata_81,
	d_writedata_22,
	readdata_22,
	readdata_71,
	readdata_61,
	readdata_20,
	d_writedata_20,
	readdata_19,
	d_writedata_19,
	src_payload7,
	src_payload8,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_411,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	out_data_buffer_313,
	out_data_buffer_314,
	out_data_buffer_302,
	out_data_buffer_303,
	out_data_buffer_292,
	out_data_buffer_293,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_data_33,
	src_payload14,
	src_payload15,
	src_data_34,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_data_35,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	av_ld_getting_data,
	src_data_51,
	src_data_71,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_28;
output 	W_alu_result_27;
output 	W_alu_result_26;
output 	W_alu_result_25;
output 	W_alu_result_24;
output 	W_alu_result_23;
output 	W_alu_result_22;
output 	W_alu_result_21;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_6;
output 	W_alu_result_7;
output 	W_alu_result_5;
output 	W_alu_result_4;
output 	W_alu_result_12;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_11;
output 	W_alu_result_2;
output 	W_alu_result_3;
input 	q_a_0;
input 	readdata_0;
input 	q_a_1;
input 	readdata_1;
input 	readdata_2;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_11;
input 	q_a_13;
input 	q_a_16;
input 	q_a_12;
input 	q_a_5;
input 	q_a_14;
input 	q_a_15;
input 	q_a_21;
input 	q_a_18;
input 	readdata_17;
input 	q_a_17;
input 	q_a_31;
input 	q_a_30;
input 	q_a_29;
input 	q_a_28;
input 	q_a_27;
input 	q_a_26;
input 	q_a_25;
input 	q_a_10;
input 	q_a_24;
input 	q_a_9;
input 	q_a_23;
input 	readdata_8;
input 	q_a_8;
input 	q_a_22;
input 	q_a_7;
input 	q_a_6;
input 	q_a_20;
input 	q_a_19;
output 	readdata_01;
output 	readdata_11;
output 	readdata_21;
output 	readdata_3;
output 	d_writedata_31;
output 	d_writedata_30;
output 	d_writedata_29;
output 	d_writedata_28;
output 	d_writedata_27;
output 	d_writedata_26;
output 	d_writedata_25;
output 	d_writedata_24;
output 	ir_out_0;
output 	ir_out_1;
output 	d_read;
output 	d_write;
output 	F_pc_26;
output 	F_pc_25;
output 	F_pc_24;
output 	F_pc_23;
output 	F_pc_22;
output 	F_pc_21;
output 	F_pc_20;
output 	F_pc_19;
output 	F_pc_18;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_5;
output 	F_pc_3;
output 	i_read;
output 	F_pc_2;
output 	F_pc_4;
output 	F_pc_9;
output 	d_writedata_0;
output 	d_byteenable_0;
output 	F_pc_0;
output 	F_pc_1;
input 	r_sync_rst;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_10;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	mem_86_0;
input 	mem_68_0;
input 	src0_valid;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	src0_valid1;
input 	src0_valid2;
input 	read_latency_shift_reg_04;
input 	mem_86_01;
input 	mem_68_01;
input 	src0_valid3;
input 	src0_valid4;
input 	WideOr1;
input 	mem_67_0;
input 	mem_67_01;
input 	mem_67_02;
input 	mem_67_03;
input 	mem_67_04;
input 	mem_67_05;
input 	mem_67_06;
input 	out_data_buffer_67;
input 	out_data_buffer_671;
input 	mem_67_07;
input 	src_payload;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	src_payload1;
input 	src_payload2;
input 	out_valid2;
input 	out_valid3;
input 	av_readdatavalid;
input 	WideOr11;
input 	local_read;
output 	hbreak_enabled;
input 	av_readdata_pre_30;
input 	src_payload3;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	out_data_buffer_0;
input 	out_data_buffer_01;
input 	av_readdata_pre_1;
input 	out_data_buffer_1;
input 	av_readdata_pre_11;
input 	out_data_buffer_11;
input 	av_readdata_pre_2;
input 	out_data_buffer_2;
input 	out_data_buffer_21;
input 	av_readdata_pre_3;
input 	readdata_31;
input 	out_data_buffer_3;
input 	out_data_buffer_31;
input 	av_readdata_pre_4;
input 	readdata_4;
input 	out_data_buffer_4;
input 	out_data_buffer_41;
output 	d_byteenable_2;
input 	mem;
input 	src_data_46;
input 	av_readdata_pre_111;
input 	out_data_buffer_111;
input 	out_data_buffer_112;
input 	av_readdata_pre_13;
input 	out_data_buffer_13;
input 	out_data_buffer_131;
input 	src_payload4;
input 	av_readdata_pre_16;
input 	out_data_buffer_16;
input 	out_data_buffer_161;
input 	av_readdata_pre_12;
input 	out_data_buffer_12;
input 	out_data_buffer_121;
input 	src_payload5;
input 	av_readdata_pre_5;
input 	out_data_buffer_5;
input 	out_data_buffer_51;
input 	out_data_buffer_14;
input 	av_readdata_pre_14;
input 	out_data_buffer_141;
input 	av_readdata_pre_15;
input 	out_data_buffer_15;
input 	out_data_buffer_151;
input 	av_readdata_pre_21;
input 	out_data_buffer_211;
input 	out_data_buffer_212;
input 	out_data_buffer_18;
input 	av_readdata_pre_18;
input 	out_data_buffer_181;
input 	av_readdata_pre_17;
input 	out_data_buffer_17;
input 	out_data_buffer_171;
input 	av_readdata_pre_31;
input 	out_data_buffer_311;
input 	out_data_buffer_312;
input 	out_data_buffer_30;
input 	av_readdata_pre_301;
input 	out_data_buffer_301;
input 	av_readdata_pre_29;
input 	out_data_buffer_29;
input 	out_data_buffer_291;
input 	out_data_buffer_28;
input 	av_readdata_pre_28;
input 	out_data_buffer_281;
input 	av_readdata_pre_27;
input 	out_data_buffer_27;
input 	out_data_buffer_271;
input 	out_data_buffer_26;
input 	av_readdata_pre_26;
input 	out_data_buffer_261;
input 	av_readdata_pre_25;
input 	out_data_buffer_25;
input 	out_data_buffer_251;
input 	out_data_buffer_10;
input 	av_readdata_pre_10;
input 	out_data_buffer_101;
input 	out_data_buffer_24;
input 	av_readdata_pre_24;
input 	out_data_buffer_241;
input 	av_readdata_pre_9;
input 	out_data_buffer_9;
input 	out_data_buffer_91;
input 	av_readdata_pre_23;
input 	out_data_buffer_23;
input 	out_data_buffer_231;
input 	out_data_buffer_8;
input 	av_readdata_pre_8;
input 	out_data_buffer_81;
input 	out_data_buffer_22;
input 	av_readdata_pre_22;
input 	out_data_buffer_221;
input 	readdata_7;
input 	out_data_buffer_7;
input 	av_readdata_pre_7;
input 	out_data_buffer_71;
input 	readdata_6;
input 	av_readdata_pre_6;
input 	out_data_buffer_6;
input 	out_data_buffer_61;
input 	av_readdata_pre_20;
input 	out_data_buffer_20;
input 	out_data_buffer_201;
input 	av_readdata_pre_19;
input 	out_data_buffer_19;
input 	out_data_buffer_191;
input 	src_payload6;
input 	src_data_0;
input 	av_readdata_9;
input 	av_readdata_8;
input 	dreg_1;
input 	r_early_rst;
output 	readdata_41;
input 	src_data_1;
input 	src_data_11;
input 	src_data_2;
input 	src_data_21;
input 	src_data_3;
input 	src_data_31;
input 	src_data_4;
input 	src_data_41;
input 	src_data_5;
input 	src_data_6;
input 	src_data_61;
input 	src_data_7;
input 	src_data_8;
input 	src_data_9;
input 	src_data_10;
input 	src_data_111;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_data_17;
output 	d_byteenable_1;
output 	d_byteenable_3;
output 	readdata_111;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
input 	out_data_buffer_282;
input 	out_data_buffer_283;
output 	readdata_211;
output 	d_writedata_21;
output 	d_writedata_18;
output 	readdata_18;
input 	out_data_buffer_272;
input 	out_data_buffer_273;
output 	readdata_171;
output 	readdata_311;
input 	out_data_buffer_262;
input 	out_data_buffer_263;
output 	readdata_30;
input 	out_data_buffer_252;
input 	out_data_buffer_253;
output 	readdata_29;
input 	out_data_buffer_242;
input 	out_data_buffer_243;
output 	readdata_28;
input 	src_data_23;
output 	readdata_27;
input 	src_data_22;
output 	readdata_26;
input 	src_data_211;
output 	readdata_25;
input 	src_data_20;
output 	readdata_10;
output 	readdata_24;
input 	src_data_19;
output 	readdata_9;
output 	d_writedata_23;
output 	readdata_23;
input 	src_data_18;
output 	readdata_81;
output 	d_writedata_22;
output 	readdata_22;
output 	readdata_71;
output 	readdata_61;
output 	readdata_20;
output 	d_writedata_20;
output 	readdata_19;
output 	d_writedata_19;
input 	src_payload7;
input 	src_payload8;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_411;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
input 	out_data_buffer_313;
input 	out_data_buffer_314;
input 	out_data_buffer_302;
input 	out_data_buffer_303;
input 	out_data_buffer_292;
input 	out_data_buffer_293;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_data_33;
input 	src_payload14;
input 	src_payload15;
input 	src_data_34;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_data_35;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
output 	av_ld_getting_data;
input 	src_data_51;
input 	src_data_71;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_final_project_soc_nios2_qsys_0_cpu cpu(
	.sr_0(sr_0),
	.W_alu_result_28(W_alu_result_28),
	.W_alu_result_27(W_alu_result_27),
	.W_alu_result_26(W_alu_result_26),
	.W_alu_result_25(W_alu_result_25),
	.W_alu_result_24(W_alu_result_24),
	.W_alu_result_23(W_alu_result_23),
	.W_alu_result_22(W_alu_result_22),
	.W_alu_result_21(W_alu_result_21),
	.W_alu_result_20(W_alu_result_20),
	.W_alu_result_19(W_alu_result_19),
	.W_alu_result_18(W_alu_result_18),
	.W_alu_result_17(W_alu_result_17),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_2(W_alu_result_2),
	.W_alu_result_3(W_alu_result_3),
	.q_a_0(q_a_0),
	.readdata_0(readdata_0),
	.q_a_1(q_a_1),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.readdata_17(readdata_17),
	.q_a_17(q_a_17),
	.q_a_31(q_a_31),
	.q_a_30(q_a_30),
	.q_a_29(q_a_29),
	.q_a_28(q_a_28),
	.q_a_27(q_a_27),
	.q_a_26(q_a_26),
	.q_a_25(q_a_25),
	.q_a_10(q_a_10),
	.q_a_24(q_a_24),
	.q_a_9(q_a_9),
	.q_a_23(q_a_23),
	.readdata_8(readdata_8),
	.q_a_8(q_a_8),
	.q_a_22(q_a_22),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.readdata_01(readdata_01),
	.readdata_11(readdata_11),
	.readdata_21(readdata_21),
	.readdata_3(readdata_3),
	.d_writedata_31(d_writedata_31),
	.d_writedata_30(d_writedata_30),
	.d_writedata_29(d_writedata_29),
	.d_writedata_28(d_writedata_28),
	.d_writedata_27(d_writedata_27),
	.d_writedata_26(d_writedata_26),
	.d_writedata_25(d_writedata_25),
	.d_writedata_24(d_writedata_24),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_read1(d_read),
	.d_write1(d_write),
	.F_pc_26(F_pc_26),
	.F_pc_25(F_pc_25),
	.F_pc_24(F_pc_24),
	.F_pc_23(F_pc_23),
	.F_pc_22(F_pc_22),
	.F_pc_21(F_pc_21),
	.F_pc_20(F_pc_20),
	.F_pc_19(F_pc_19),
	.F_pc_18(F_pc_18),
	.F_pc_17(F_pc_17),
	.F_pc_16(F_pc_16),
	.F_pc_15(F_pc_15),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.F_pc_10(F_pc_10),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_3(F_pc_3),
	.i_read1(i_read),
	.F_pc_2(F_pc_2),
	.F_pc_4(F_pc_4),
	.F_pc_9(F_pc_9),
	.d_writedata_0(d_writedata_0),
	.d_byteenable_0(d_byteenable_0),
	.F_pc_0(F_pc_0),
	.F_pc_1(F_pc_1),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.d_writedata_8(d_writedata_8),
	.d_writedata_9(d_writedata_9),
	.d_writedata_10(d_writedata_10),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_17(d_writedata_17),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.mem_86_0(mem_86_0),
	.mem_68_0(mem_68_0),
	.src0_valid(src0_valid),
	.out_valid(out_valid),
	.out_data_toggle_flopped(out_data_toggle_flopped),
	.dreg_0(dreg_0),
	.out_valid1(out_valid1),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.read_latency_shift_reg_03(read_latency_shift_reg_03),
	.src0_valid1(src0_valid1),
	.src0_valid2(src0_valid2),
	.read_latency_shift_reg_04(read_latency_shift_reg_04),
	.mem_86_01(mem_86_01),
	.mem_68_01(mem_68_01),
	.src0_valid3(src0_valid3),
	.src0_valid4(src0_valid4),
	.WideOr1(WideOr1),
	.mem_67_0(mem_67_0),
	.mem_67_01(mem_67_01),
	.mem_67_02(mem_67_02),
	.mem_67_03(mem_67_03),
	.mem_67_04(mem_67_04),
	.mem_67_05(mem_67_05),
	.mem_67_06(mem_67_06),
	.out_data_buffer_67(out_data_buffer_67),
	.out_data_buffer_671(out_data_buffer_671),
	.mem_67_07(mem_67_07),
	.src_payload(src_payload),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.av_waitrequest(av_waitrequest),
	.src1_valid(src1_valid),
	.src1_valid1(src1_valid1),
	.src1_valid2(src1_valid2),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.out_valid2(out_valid2),
	.out_valid3(out_valid3),
	.av_readdatavalid(av_readdatavalid),
	.WideOr11(WideOr11),
	.local_read(local_read),
	.hbreak_enabled1(hbreak_enabled),
	.av_readdata_pre_30(av_readdata_pre_30),
	.src_payload3(src_payload3),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_01(av_readdata_pre_01),
	.out_data_buffer_0(out_data_buffer_0),
	.out_data_buffer_01(out_data_buffer_01),
	.av_readdata_pre_1(av_readdata_pre_1),
	.out_data_buffer_1(out_data_buffer_1),
	.av_readdata_pre_11(av_readdata_pre_11),
	.out_data_buffer_11(out_data_buffer_11),
	.av_readdata_pre_2(av_readdata_pre_2),
	.out_data_buffer_2(out_data_buffer_2),
	.out_data_buffer_21(out_data_buffer_21),
	.av_readdata_pre_3(av_readdata_pre_3),
	.readdata_31(readdata_31),
	.out_data_buffer_3(out_data_buffer_3),
	.out_data_buffer_31(out_data_buffer_31),
	.av_readdata_pre_4(av_readdata_pre_4),
	.readdata_4(readdata_4),
	.out_data_buffer_4(out_data_buffer_4),
	.out_data_buffer_41(out_data_buffer_41),
	.d_byteenable_2(d_byteenable_2),
	.mem(mem),
	.src_data_46(src_data_46),
	.av_readdata_pre_111(av_readdata_pre_111),
	.out_data_buffer_111(out_data_buffer_111),
	.out_data_buffer_112(out_data_buffer_112),
	.av_readdata_pre_13(av_readdata_pre_13),
	.out_data_buffer_13(out_data_buffer_13),
	.out_data_buffer_131(out_data_buffer_131),
	.src_payload4(src_payload4),
	.av_readdata_pre_16(av_readdata_pre_16),
	.out_data_buffer_16(out_data_buffer_16),
	.out_data_buffer_161(out_data_buffer_161),
	.av_readdata_pre_12(av_readdata_pre_12),
	.out_data_buffer_12(out_data_buffer_12),
	.out_data_buffer_121(out_data_buffer_121),
	.src_payload5(src_payload5),
	.av_readdata_pre_5(av_readdata_pre_5),
	.out_data_buffer_5(out_data_buffer_5),
	.out_data_buffer_51(out_data_buffer_51),
	.out_data_buffer_14(out_data_buffer_14),
	.av_readdata_pre_14(av_readdata_pre_14),
	.out_data_buffer_141(out_data_buffer_141),
	.av_readdata_pre_15(av_readdata_pre_15),
	.out_data_buffer_15(out_data_buffer_15),
	.out_data_buffer_151(out_data_buffer_151),
	.av_readdata_pre_21(av_readdata_pre_21),
	.out_data_buffer_211(out_data_buffer_211),
	.out_data_buffer_212(out_data_buffer_212),
	.out_data_buffer_18(out_data_buffer_18),
	.av_readdata_pre_18(av_readdata_pre_18),
	.out_data_buffer_181(out_data_buffer_181),
	.av_readdata_pre_17(av_readdata_pre_17),
	.out_data_buffer_17(out_data_buffer_17),
	.out_data_buffer_171(out_data_buffer_171),
	.av_readdata_pre_31(av_readdata_pre_31),
	.out_data_buffer_311(out_data_buffer_311),
	.out_data_buffer_312(out_data_buffer_312),
	.out_data_buffer_30(out_data_buffer_30),
	.av_readdata_pre_301(av_readdata_pre_301),
	.out_data_buffer_301(out_data_buffer_301),
	.av_readdata_pre_29(av_readdata_pre_29),
	.out_data_buffer_29(out_data_buffer_29),
	.out_data_buffer_291(out_data_buffer_291),
	.out_data_buffer_28(out_data_buffer_28),
	.av_readdata_pre_28(av_readdata_pre_28),
	.out_data_buffer_281(out_data_buffer_281),
	.av_readdata_pre_27(av_readdata_pre_27),
	.out_data_buffer_27(out_data_buffer_27),
	.out_data_buffer_271(out_data_buffer_271),
	.out_data_buffer_26(out_data_buffer_26),
	.av_readdata_pre_26(av_readdata_pre_26),
	.out_data_buffer_261(out_data_buffer_261),
	.av_readdata_pre_25(av_readdata_pre_25),
	.out_data_buffer_25(out_data_buffer_25),
	.out_data_buffer_251(out_data_buffer_251),
	.out_data_buffer_10(out_data_buffer_10),
	.av_readdata_pre_10(av_readdata_pre_10),
	.out_data_buffer_101(out_data_buffer_101),
	.out_data_buffer_24(out_data_buffer_24),
	.av_readdata_pre_24(av_readdata_pre_24),
	.out_data_buffer_241(out_data_buffer_241),
	.av_readdata_pre_9(av_readdata_pre_9),
	.out_data_buffer_9(out_data_buffer_9),
	.out_data_buffer_91(out_data_buffer_91),
	.av_readdata_pre_23(av_readdata_pre_23),
	.out_data_buffer_23(out_data_buffer_23),
	.out_data_buffer_231(out_data_buffer_231),
	.out_data_buffer_8(out_data_buffer_8),
	.av_readdata_pre_8(av_readdata_pre_8),
	.out_data_buffer_81(out_data_buffer_81),
	.out_data_buffer_22(out_data_buffer_22),
	.av_readdata_pre_22(av_readdata_pre_22),
	.out_data_buffer_221(out_data_buffer_221),
	.readdata_7(readdata_7),
	.out_data_buffer_7(out_data_buffer_7),
	.av_readdata_pre_7(av_readdata_pre_7),
	.out_data_buffer_71(out_data_buffer_71),
	.readdata_6(readdata_6),
	.av_readdata_pre_6(av_readdata_pre_6),
	.out_data_buffer_6(out_data_buffer_6),
	.out_data_buffer_61(out_data_buffer_61),
	.av_readdata_pre_20(av_readdata_pre_20),
	.out_data_buffer_20(out_data_buffer_20),
	.out_data_buffer_201(out_data_buffer_201),
	.av_readdata_pre_19(av_readdata_pre_19),
	.out_data_buffer_19(out_data_buffer_19),
	.out_data_buffer_191(out_data_buffer_191),
	.src_payload6(src_payload6),
	.src_data_0(src_data_0),
	.av_readdata_9(av_readdata_9),
	.av_readdata_8(av_readdata_8),
	.dreg_1(dreg_1),
	.r_early_rst(r_early_rst),
	.readdata_41(readdata_41),
	.src_data_1(src_data_1),
	.src_data_11(src_data_11),
	.src_data_2(src_data_2),
	.src_data_21(src_data_21),
	.src_data_3(src_data_3),
	.src_data_31(src_data_31),
	.src_data_4(src_data_4),
	.src_data_41(src_data_41),
	.src_data_5(src_data_5),
	.src_data_6(src_data_6),
	.src_data_61(src_data_61),
	.src_data_7(src_data_7),
	.src_data_8(src_data_8),
	.src_data_9(src_data_9),
	.src_data_10(src_data_10),
	.src_data_111(src_data_111),
	.src_data_12(src_data_12),
	.src_data_13(src_data_13),
	.src_data_14(src_data_14),
	.src_data_15(src_data_15),
	.src_data_16(src_data_16),
	.src_data_17(src_data_17),
	.d_byteenable_1(d_byteenable_1),
	.d_byteenable_3(d_byteenable_3),
	.readdata_111(readdata_111),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_5(readdata_5),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.out_data_buffer_282(out_data_buffer_282),
	.out_data_buffer_283(out_data_buffer_283),
	.readdata_211(readdata_211),
	.d_writedata_21(d_writedata_21),
	.d_writedata_18(d_writedata_18),
	.readdata_18(readdata_18),
	.out_data_buffer_272(out_data_buffer_272),
	.out_data_buffer_273(out_data_buffer_273),
	.readdata_171(readdata_171),
	.readdata_311(readdata_311),
	.out_data_buffer_262(out_data_buffer_262),
	.out_data_buffer_263(out_data_buffer_263),
	.readdata_30(readdata_30),
	.out_data_buffer_252(out_data_buffer_252),
	.out_data_buffer_253(out_data_buffer_253),
	.readdata_29(readdata_29),
	.out_data_buffer_242(out_data_buffer_242),
	.out_data_buffer_243(out_data_buffer_243),
	.readdata_28(readdata_28),
	.src_data_23(src_data_23),
	.readdata_27(readdata_27),
	.src_data_22(src_data_22),
	.readdata_26(readdata_26),
	.src_data_211(src_data_211),
	.readdata_25(readdata_25),
	.src_data_20(src_data_20),
	.readdata_10(readdata_10),
	.readdata_24(readdata_24),
	.src_data_19(src_data_19),
	.readdata_9(readdata_9),
	.d_writedata_23(d_writedata_23),
	.readdata_23(readdata_23),
	.src_data_18(src_data_18),
	.readdata_81(readdata_81),
	.d_writedata_22(d_writedata_22),
	.readdata_22(readdata_22),
	.readdata_71(readdata_71),
	.readdata_61(readdata_61),
	.readdata_20(readdata_20),
	.d_writedata_20(d_writedata_20),
	.readdata_19(readdata_19),
	.d_writedata_19(d_writedata_19),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_411(src_data_411),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.out_data_buffer_313(out_data_buffer_313),
	.out_data_buffer_314(out_data_buffer_314),
	.out_data_buffer_302(out_data_buffer_302),
	.out_data_buffer_303(out_data_buffer_303),
	.out_data_buffer_292(out_data_buffer_292),
	.out_data_buffer_293(out_data_buffer_293),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_data_33(src_data_33),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_data_34(src_data_34),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_data_35(src_data_35),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.src_payload33(src_payload33),
	.src_payload34(src_payload34),
	.src_payload35(src_payload35),
	.src_payload36(src_payload36),
	.src_payload37(src_payload37),
	.src_payload38(src_payload38),
	.src_payload39(src_payload39),
	.av_ld_getting_data(av_ld_getting_data),
	.src_data_51(src_data_51),
	.src_data_71(src_data_71),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu (
	sr_0,
	W_alu_result_28,
	W_alu_result_27,
	W_alu_result_26,
	W_alu_result_25,
	W_alu_result_24,
	W_alu_result_23,
	W_alu_result_22,
	W_alu_result_21,
	W_alu_result_20,
	W_alu_result_19,
	W_alu_result_18,
	W_alu_result_17,
	W_alu_result_16,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_6,
	W_alu_result_7,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_12,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_11,
	W_alu_result_2,
	W_alu_result_3,
	q_a_0,
	readdata_0,
	q_a_1,
	readdata_1,
	readdata_2,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	readdata_17,
	q_a_17,
	q_a_31,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_10,
	q_a_24,
	q_a_9,
	q_a_23,
	readdata_8,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	readdata_01,
	readdata_11,
	readdata_21,
	readdata_3,
	d_writedata_31,
	d_writedata_30,
	d_writedata_29,
	d_writedata_28,
	d_writedata_27,
	d_writedata_26,
	d_writedata_25,
	d_writedata_24,
	ir_out_0,
	ir_out_1,
	d_read1,
	d_write1,
	F_pc_26,
	F_pc_25,
	F_pc_24,
	F_pc_23,
	F_pc_22,
	F_pc_21,
	F_pc_20,
	F_pc_19,
	F_pc_18,
	F_pc_17,
	F_pc_16,
	F_pc_15,
	F_pc_14,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	F_pc_10,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_3,
	i_read1,
	F_pc_2,
	F_pc_4,
	F_pc_9,
	d_writedata_0,
	d_byteenable_0,
	F_pc_0,
	F_pc_1,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	d_writedata_8,
	d_writedata_9,
	d_writedata_10,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_17,
	read_latency_shift_reg_0,
	read_latency_shift_reg_01,
	mem_86_0,
	mem_68_0,
	src0_valid,
	out_valid,
	out_data_toggle_flopped,
	dreg_0,
	out_valid1,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	src0_valid1,
	src0_valid2,
	read_latency_shift_reg_04,
	mem_86_01,
	mem_68_01,
	src0_valid3,
	src0_valid4,
	WideOr1,
	mem_67_0,
	mem_67_01,
	mem_67_02,
	mem_67_03,
	mem_67_04,
	mem_67_05,
	mem_67_06,
	out_data_buffer_67,
	out_data_buffer_671,
	mem_67_07,
	src_payload,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	src1_valid,
	src1_valid1,
	src1_valid2,
	src_payload1,
	src_payload2,
	out_valid2,
	out_valid3,
	av_readdatavalid,
	WideOr11,
	local_read,
	hbreak_enabled1,
	av_readdata_pre_30,
	src_payload3,
	av_readdata_pre_0,
	av_readdata_pre_01,
	out_data_buffer_0,
	out_data_buffer_01,
	av_readdata_pre_1,
	out_data_buffer_1,
	av_readdata_pre_11,
	out_data_buffer_11,
	av_readdata_pre_2,
	out_data_buffer_2,
	out_data_buffer_21,
	av_readdata_pre_3,
	readdata_31,
	out_data_buffer_3,
	out_data_buffer_31,
	av_readdata_pre_4,
	readdata_4,
	out_data_buffer_4,
	out_data_buffer_41,
	d_byteenable_2,
	mem,
	src_data_46,
	av_readdata_pre_111,
	out_data_buffer_111,
	out_data_buffer_112,
	av_readdata_pre_13,
	out_data_buffer_13,
	out_data_buffer_131,
	src_payload4,
	av_readdata_pre_16,
	out_data_buffer_16,
	out_data_buffer_161,
	av_readdata_pre_12,
	out_data_buffer_12,
	out_data_buffer_121,
	src_payload5,
	av_readdata_pre_5,
	out_data_buffer_5,
	out_data_buffer_51,
	out_data_buffer_14,
	av_readdata_pre_14,
	out_data_buffer_141,
	av_readdata_pre_15,
	out_data_buffer_15,
	out_data_buffer_151,
	av_readdata_pre_21,
	out_data_buffer_211,
	out_data_buffer_212,
	out_data_buffer_18,
	av_readdata_pre_18,
	out_data_buffer_181,
	av_readdata_pre_17,
	out_data_buffer_17,
	out_data_buffer_171,
	av_readdata_pre_31,
	out_data_buffer_311,
	out_data_buffer_312,
	out_data_buffer_30,
	av_readdata_pre_301,
	out_data_buffer_301,
	av_readdata_pre_29,
	out_data_buffer_29,
	out_data_buffer_291,
	out_data_buffer_28,
	av_readdata_pre_28,
	out_data_buffer_281,
	av_readdata_pre_27,
	out_data_buffer_27,
	out_data_buffer_271,
	out_data_buffer_26,
	av_readdata_pre_26,
	out_data_buffer_261,
	av_readdata_pre_25,
	out_data_buffer_25,
	out_data_buffer_251,
	out_data_buffer_10,
	av_readdata_pre_10,
	out_data_buffer_101,
	out_data_buffer_24,
	av_readdata_pre_24,
	out_data_buffer_241,
	av_readdata_pre_9,
	out_data_buffer_9,
	out_data_buffer_91,
	av_readdata_pre_23,
	out_data_buffer_23,
	out_data_buffer_231,
	out_data_buffer_8,
	av_readdata_pre_8,
	out_data_buffer_81,
	out_data_buffer_22,
	av_readdata_pre_22,
	out_data_buffer_221,
	readdata_7,
	out_data_buffer_7,
	av_readdata_pre_7,
	out_data_buffer_71,
	readdata_6,
	av_readdata_pre_6,
	out_data_buffer_6,
	out_data_buffer_61,
	av_readdata_pre_20,
	out_data_buffer_20,
	out_data_buffer_201,
	av_readdata_pre_19,
	out_data_buffer_19,
	out_data_buffer_191,
	src_payload6,
	src_data_0,
	av_readdata_9,
	av_readdata_8,
	dreg_1,
	r_early_rst,
	readdata_41,
	src_data_1,
	src_data_11,
	src_data_2,
	src_data_21,
	src_data_3,
	src_data_31,
	src_data_4,
	src_data_41,
	src_data_5,
	src_data_6,
	src_data_61,
	src_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_111,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	d_byteenable_1,
	d_byteenable_3,
	readdata_111,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	out_data_buffer_282,
	out_data_buffer_283,
	readdata_211,
	d_writedata_21,
	d_writedata_18,
	readdata_18,
	out_data_buffer_272,
	out_data_buffer_273,
	readdata_171,
	readdata_311,
	out_data_buffer_262,
	out_data_buffer_263,
	readdata_30,
	out_data_buffer_252,
	out_data_buffer_253,
	readdata_29,
	out_data_buffer_242,
	out_data_buffer_243,
	readdata_28,
	src_data_23,
	readdata_27,
	src_data_22,
	readdata_26,
	src_data_211,
	readdata_25,
	src_data_20,
	readdata_10,
	readdata_24,
	src_data_19,
	readdata_9,
	d_writedata_23,
	readdata_23,
	src_data_18,
	readdata_81,
	d_writedata_22,
	readdata_22,
	readdata_71,
	readdata_61,
	readdata_20,
	d_writedata_20,
	readdata_19,
	d_writedata_19,
	src_payload7,
	src_payload8,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_411,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	out_data_buffer_313,
	out_data_buffer_314,
	out_data_buffer_302,
	out_data_buffer_303,
	out_data_buffer_292,
	out_data_buffer_293,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_data_33,
	src_payload14,
	src_payload15,
	src_data_34,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_data_35,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	av_ld_getting_data,
	src_data_51,
	src_data_71,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_28;
output 	W_alu_result_27;
output 	W_alu_result_26;
output 	W_alu_result_25;
output 	W_alu_result_24;
output 	W_alu_result_23;
output 	W_alu_result_22;
output 	W_alu_result_21;
output 	W_alu_result_20;
output 	W_alu_result_19;
output 	W_alu_result_18;
output 	W_alu_result_17;
output 	W_alu_result_16;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_6;
output 	W_alu_result_7;
output 	W_alu_result_5;
output 	W_alu_result_4;
output 	W_alu_result_12;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_11;
output 	W_alu_result_2;
output 	W_alu_result_3;
input 	q_a_0;
input 	readdata_0;
input 	q_a_1;
input 	readdata_1;
input 	readdata_2;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_11;
input 	q_a_13;
input 	q_a_16;
input 	q_a_12;
input 	q_a_5;
input 	q_a_14;
input 	q_a_15;
input 	q_a_21;
input 	q_a_18;
input 	readdata_17;
input 	q_a_17;
input 	q_a_31;
input 	q_a_30;
input 	q_a_29;
input 	q_a_28;
input 	q_a_27;
input 	q_a_26;
input 	q_a_25;
input 	q_a_10;
input 	q_a_24;
input 	q_a_9;
input 	q_a_23;
input 	readdata_8;
input 	q_a_8;
input 	q_a_22;
input 	q_a_7;
input 	q_a_6;
input 	q_a_20;
input 	q_a_19;
output 	readdata_01;
output 	readdata_11;
output 	readdata_21;
output 	readdata_3;
output 	d_writedata_31;
output 	d_writedata_30;
output 	d_writedata_29;
output 	d_writedata_28;
output 	d_writedata_27;
output 	d_writedata_26;
output 	d_writedata_25;
output 	d_writedata_24;
output 	ir_out_0;
output 	ir_out_1;
output 	d_read1;
output 	d_write1;
output 	F_pc_26;
output 	F_pc_25;
output 	F_pc_24;
output 	F_pc_23;
output 	F_pc_22;
output 	F_pc_21;
output 	F_pc_20;
output 	F_pc_19;
output 	F_pc_18;
output 	F_pc_17;
output 	F_pc_16;
output 	F_pc_15;
output 	F_pc_14;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	F_pc_10;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_5;
output 	F_pc_3;
output 	i_read1;
output 	F_pc_2;
output 	F_pc_4;
output 	F_pc_9;
output 	d_writedata_0;
output 	d_byteenable_0;
output 	F_pc_0;
output 	F_pc_1;
input 	r_sync_rst;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
output 	d_writedata_8;
output 	d_writedata_9;
output 	d_writedata_10;
output 	d_writedata_11;
output 	d_writedata_12;
output 	d_writedata_13;
output 	d_writedata_14;
output 	d_writedata_15;
output 	d_writedata_16;
output 	d_writedata_17;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_01;
input 	mem_86_0;
input 	mem_68_0;
input 	src0_valid;
input 	out_valid;
input 	out_data_toggle_flopped;
input 	dreg_0;
input 	out_valid1;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	src0_valid1;
input 	src0_valid2;
input 	read_latency_shift_reg_04;
input 	mem_86_01;
input 	mem_68_01;
input 	src0_valid3;
input 	src0_valid4;
input 	WideOr1;
input 	mem_67_0;
input 	mem_67_01;
input 	mem_67_02;
input 	mem_67_03;
input 	mem_67_04;
input 	mem_67_05;
input 	mem_67_06;
input 	out_data_buffer_67;
input 	out_data_buffer_671;
input 	mem_67_07;
input 	src_payload;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
input 	src1_valid;
input 	src1_valid1;
input 	src1_valid2;
input 	src_payload1;
input 	src_payload2;
input 	out_valid2;
input 	out_valid3;
input 	av_readdatavalid;
input 	WideOr11;
input 	local_read;
output 	hbreak_enabled1;
input 	av_readdata_pre_30;
input 	src_payload3;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	out_data_buffer_0;
input 	out_data_buffer_01;
input 	av_readdata_pre_1;
input 	out_data_buffer_1;
input 	av_readdata_pre_11;
input 	out_data_buffer_11;
input 	av_readdata_pre_2;
input 	out_data_buffer_2;
input 	out_data_buffer_21;
input 	av_readdata_pre_3;
input 	readdata_31;
input 	out_data_buffer_3;
input 	out_data_buffer_31;
input 	av_readdata_pre_4;
input 	readdata_4;
input 	out_data_buffer_4;
input 	out_data_buffer_41;
output 	d_byteenable_2;
input 	mem;
input 	src_data_46;
input 	av_readdata_pre_111;
input 	out_data_buffer_111;
input 	out_data_buffer_112;
input 	av_readdata_pre_13;
input 	out_data_buffer_13;
input 	out_data_buffer_131;
input 	src_payload4;
input 	av_readdata_pre_16;
input 	out_data_buffer_16;
input 	out_data_buffer_161;
input 	av_readdata_pre_12;
input 	out_data_buffer_12;
input 	out_data_buffer_121;
input 	src_payload5;
input 	av_readdata_pre_5;
input 	out_data_buffer_5;
input 	out_data_buffer_51;
input 	out_data_buffer_14;
input 	av_readdata_pre_14;
input 	out_data_buffer_141;
input 	av_readdata_pre_15;
input 	out_data_buffer_15;
input 	out_data_buffer_151;
input 	av_readdata_pre_21;
input 	out_data_buffer_211;
input 	out_data_buffer_212;
input 	out_data_buffer_18;
input 	av_readdata_pre_18;
input 	out_data_buffer_181;
input 	av_readdata_pre_17;
input 	out_data_buffer_17;
input 	out_data_buffer_171;
input 	av_readdata_pre_31;
input 	out_data_buffer_311;
input 	out_data_buffer_312;
input 	out_data_buffer_30;
input 	av_readdata_pre_301;
input 	out_data_buffer_301;
input 	av_readdata_pre_29;
input 	out_data_buffer_29;
input 	out_data_buffer_291;
input 	out_data_buffer_28;
input 	av_readdata_pre_28;
input 	out_data_buffer_281;
input 	av_readdata_pre_27;
input 	out_data_buffer_27;
input 	out_data_buffer_271;
input 	out_data_buffer_26;
input 	av_readdata_pre_26;
input 	out_data_buffer_261;
input 	av_readdata_pre_25;
input 	out_data_buffer_25;
input 	out_data_buffer_251;
input 	out_data_buffer_10;
input 	av_readdata_pre_10;
input 	out_data_buffer_101;
input 	out_data_buffer_24;
input 	av_readdata_pre_24;
input 	out_data_buffer_241;
input 	av_readdata_pre_9;
input 	out_data_buffer_9;
input 	out_data_buffer_91;
input 	av_readdata_pre_23;
input 	out_data_buffer_23;
input 	out_data_buffer_231;
input 	out_data_buffer_8;
input 	av_readdata_pre_8;
input 	out_data_buffer_81;
input 	out_data_buffer_22;
input 	av_readdata_pre_22;
input 	out_data_buffer_221;
input 	readdata_7;
input 	out_data_buffer_7;
input 	av_readdata_pre_7;
input 	out_data_buffer_71;
input 	readdata_6;
input 	av_readdata_pre_6;
input 	out_data_buffer_6;
input 	out_data_buffer_61;
input 	av_readdata_pre_20;
input 	out_data_buffer_20;
input 	out_data_buffer_201;
input 	av_readdata_pre_19;
input 	out_data_buffer_19;
input 	out_data_buffer_191;
input 	src_payload6;
input 	src_data_0;
input 	av_readdata_9;
input 	av_readdata_8;
input 	dreg_1;
input 	r_early_rst;
output 	readdata_41;
input 	src_data_1;
input 	src_data_11;
input 	src_data_2;
input 	src_data_21;
input 	src_data_3;
input 	src_data_31;
input 	src_data_4;
input 	src_data_41;
input 	src_data_5;
input 	src_data_6;
input 	src_data_61;
input 	src_data_7;
input 	src_data_8;
input 	src_data_9;
input 	src_data_10;
input 	src_data_111;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_data_17;
output 	d_byteenable_1;
output 	d_byteenable_3;
output 	readdata_111;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
input 	out_data_buffer_282;
input 	out_data_buffer_283;
output 	readdata_211;
output 	d_writedata_21;
output 	d_writedata_18;
output 	readdata_18;
input 	out_data_buffer_272;
input 	out_data_buffer_273;
output 	readdata_171;
output 	readdata_311;
input 	out_data_buffer_262;
input 	out_data_buffer_263;
output 	readdata_30;
input 	out_data_buffer_252;
input 	out_data_buffer_253;
output 	readdata_29;
input 	out_data_buffer_242;
input 	out_data_buffer_243;
output 	readdata_28;
input 	src_data_23;
output 	readdata_27;
input 	src_data_22;
output 	readdata_26;
input 	src_data_211;
output 	readdata_25;
input 	src_data_20;
output 	readdata_10;
output 	readdata_24;
input 	src_data_19;
output 	readdata_9;
output 	d_writedata_23;
output 	readdata_23;
input 	src_data_18;
output 	readdata_81;
output 	d_writedata_22;
output 	readdata_22;
output 	readdata_71;
output 	readdata_61;
output 	readdata_20;
output 	d_writedata_20;
output 	readdata_19;
output 	d_writedata_19;
input 	src_payload7;
input 	src_payload8;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_411;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
input 	out_data_buffer_313;
input 	out_data_buffer_314;
input 	out_data_buffer_302;
input 	out_data_buffer_303;
input 	out_data_buffer_292;
input 	out_data_buffer_293;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_data_33;
input 	src_payload14;
input 	src_payload15;
input 	src_data_34;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_data_35;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
output 	av_ld_getting_data;
input 	src_data_51;
input 	src_data_71;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \Add1~92_combout ;
wire \Add1~94_combout ;
wire \Add1~96_combout ;
wire \W_alu_result[0]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|jtag_break~q ;
wire \W_alu_result[1]~q ;
wire \av_ld_byte1_data[0]~q ;
wire \av_ld_byte1_data[1]~q ;
wire \av_ld_byte1_data[2]~q ;
wire \av_ld_byte1_data[3]~q ;
wire \av_ld_byte1_data[4]~q ;
wire \av_ld_byte1_data[5]~q ;
wire \av_ld_byte1_data[6]~q ;
wire \av_ld_byte1_data[7]~q ;
wire \av_ld_byte2_data[0]~q ;
wire \av_ld_byte2_data[1]~q ;
wire \av_ld_byte2_data[7]~q ;
wire \av_ld_byte2_data[6]~q ;
wire \av_ld_byte2_data[5]~q ;
wire \av_ld_byte2_data[4]~q ;
wire \av_ld_byte2_data[3]~q ;
wire \av_ld_byte2_data[2]~q ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \W_alu_result[0]~27_combout ;
wire \W_alu_result[1]~28_combout ;
wire \av_ld_byte1_data[0]~0_combout ;
wire \av_ld_byte1_data[1]~1_combout ;
wire \av_ld_byte1_data[2]~2_combout ;
wire \av_ld_byte1_data[3]~3_combout ;
wire \av_ld_byte1_data[4]~4_combout ;
wire \av_ld_byte1_data[5]~5_combout ;
wire \av_ld_byte1_data[6]~6_combout ;
wire \av_ld_byte1_data[7]~7_combout ;
wire \av_ld_byte2_data[0]~0_combout ;
wire \av_ld_byte2_data[1]~1_combout ;
wire \av_ld_byte2_data[7]~2_combout ;
wire \av_ld_byte2_data[6]~3_combout ;
wire \av_ld_byte2_data[5]~4_combout ;
wire \av_ld_byte2_data[4]~5_combout ;
wire \av_ld_byte2_data[3]~6_combout ;
wire \av_ld_byte2_data[2]~7_combout ;
wire \W_alu_result[31]~q ;
wire \W_alu_result[30]~q ;
wire \W_alu_result[29]~q ;
wire \W_alu_result[31]~29_combout ;
wire \W_alu_result[30]~30_combout ;
wire \W_alu_result[29]~31_combout ;
wire \D_ctrl_ld_signed~1_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \av_ld_byte0_data[0]~q ;
wire \W_rf_wr_data[0]~0_combout ;
wire \W_control_rd_data[0]~q ;
wire \W_rf_wr_data[0]~1_combout ;
wire \W_rf_wr_data[0]~2_combout ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \av_ld_byte0_data[1]~q ;
wire \W_control_rd_data[1]~q ;
wire \W_rf_wr_data[1]~3_combout ;
wire \W_rf_wr_data[1]~4_combout ;
wire \av_ld_byte0_data[2]~q ;
wire \W_rf_wr_data[2]~5_combout ;
wire \av_ld_byte0_data[3]~q ;
wire \W_rf_wr_data[3]~6_combout ;
wire \av_ld_byte0_data[4]~q ;
wire \W_rf_wr_data[4]~7_combout ;
wire \av_ld_byte0_data[5]~q ;
wire \W_rf_wr_data[5]~8_combout ;
wire \av_ld_byte0_data[6]~q ;
wire \W_rf_wr_data[6]~9_combout ;
wire \av_ld_byte0_data[7]~q ;
wire \W_rf_wr_data[7]~10_combout ;
wire \W_rf_wr_data[8]~11_combout ;
wire \W_rf_wr_data[9]~12_combout ;
wire \W_rf_wr_data[10]~13_combout ;
wire \W_rf_wr_data[11]~14_combout ;
wire \W_rf_wr_data[12]~15_combout ;
wire \W_rf_wr_data[13]~16_combout ;
wire \W_rf_wr_data[14]~17_combout ;
wire \W_rf_wr_data[15]~18_combout ;
wire \W_rf_wr_data[16]~19_combout ;
wire \W_rf_wr_data[17]~20_combout ;
wire \av_ld_byte3_data[4]~q ;
wire \W_rf_wr_data[28]~21_combout ;
wire \av_ld_byte3_data[3]~q ;
wire \W_rf_wr_data[27]~22_combout ;
wire \av_ld_byte3_data[2]~q ;
wire \W_rf_wr_data[26]~23_combout ;
wire \av_ld_byte3_data[1]~q ;
wire \W_rf_wr_data[25]~24_combout ;
wire \av_ld_byte3_data[0]~q ;
wire \W_rf_wr_data[24]~25_combout ;
wire \W_rf_wr_data[23]~26_combout ;
wire \W_rf_wr_data[22]~27_combout ;
wire \W_rf_wr_data[21]~28_combout ;
wire \W_rf_wr_data[20]~29_combout ;
wire \W_rf_wr_data[19]~30_combout ;
wire \W_rf_wr_data[18]~31_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~1_combout ;
wire \Equal0~17_combout ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_dst_regnum[4]~5_combout ;
wire \D_dst_regnum[4]~6_combout ;
wire \D_dst_regnum[4]~7_combout ;
wire \D_dst_regnum[4]~8_combout ;
wire \D_dst_regnum[4]~9_combout ;
wire \D_dst_regnum[0]~10_combout ;
wire \D_dst_regnum[3]~11_combout ;
wire \D_dst_regnum[2]~12_combout ;
wire \Equal0~18_combout ;
wire \D_dst_regnum[1]~13_combout ;
wire \D_dst_regnum[1]~14_combout ;
wire \D_wr_dst_reg~2_combout ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_rshift8~1_combout ;
wire \av_ld_byte0_data[1]~0_combout ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_control_rd_data[0]~1_combout ;
wire \E_control_rd_data[0]~2_combout ;
wire \E_control_rd_data[0]~3_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[1]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \av_ld_byte0_data_nxt[1]~2_combout ;
wire \E_control_rd_data[1]~4_combout ;
wire \E_control_rd_data[1]~5_combout ;
wire \av_ld_byte0_data_nxt[2]~3_combout ;
wire \av_ld_byte0_data_nxt[3]~4_combout ;
wire \av_ld_byte0_data_nxt[4]~5_combout ;
wire \av_ld_byte0_data_nxt[5]~6_combout ;
wire \av_ld_byte0_data_nxt[6]~7_combout ;
wire \av_ld_byte0_data_nxt[7]~8_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \av_ld_byte3_data_nxt~0_combout ;
wire \av_ld_byte3_data_nxt~1_combout ;
wire \av_ld_byte3_data_nxt~2_combout ;
wire \av_ld_byte3_data_nxt~3_combout ;
wire \av_ld_byte3_data_nxt~4_combout ;
wire \av_ld_byte3_data_nxt~5_combout ;
wire \av_ld_byte3_data_nxt~6_combout ;
wire \av_ld_byte3_data_nxt~7_combout ;
wire \av_ld_byte3_data_nxt~8_combout ;
wire \av_ld_byte3_data_nxt~9_combout ;
wire \av_ld_byte3_data_nxt~10_combout ;
wire \av_ld_byte3_data_nxt~11_combout ;
wire \av_ld_byte3_data_nxt~12_combout ;
wire \av_ld_byte3_data_nxt~13_combout ;
wire \av_ld_byte3_data_nxt~14_combout ;
wire \av_ld_byte3_data_nxt~15_combout ;
wire \av_ld_byte3_data_nxt~16_combout ;
wire \av_ld_byte3_data_nxt~17_combout ;
wire \av_ld_byte3_data[7]~q ;
wire \av_ld_byte3_data[6]~q ;
wire \av_ld_byte3_data[5]~q ;
wire \W_rf_wr_data[31]~32_combout ;
wire \W_rf_wr_data[30]~33_combout ;
wire \W_rf_wr_data[29]~34_combout ;
wire \av_ld_byte3_data_nxt~18_combout ;
wire \av_ld_byte3_data_nxt~19_combout ;
wire \av_ld_byte3_data_nxt~20_combout ;
wire \av_ld_byte3_data_nxt~21_combout ;
wire \av_ld_byte3_data_nxt~22_combout ;
wire \av_ld_byte3_data_nxt~23_combout ;
wire \av_ld_byte3_data_nxt~24_combout ;
wire \av_ld_byte3_data_nxt~25_combout ;
wire \av_ld_byte3_data_nxt~26_combout ;
wire \av_ld_byte3_data_nxt~27_combout ;
wire \av_ld_byte0_data_nxt[0]~9_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \av_ld_getting_data~2_combout ;
wire \av_ld_getting_data~3_combout ;
wire \av_ld_getting_data~4_combout ;
wire \av_ld_getting_data~5_combout ;
wire \av_ld_getting_data~6_combout ;
wire \av_ld_getting_data~7_combout ;
wire \av_ld_getting_data~8_combout ;
wire \E_new_inst~q ;
wire \F_iw[2]~13_combout ;
wire \F_iw[2]~14_combout ;
wire \F_iw[2]~15_combout ;
wire \F_iw[2]~16_combout ;
wire \D_iw[2]~q ;
wire \F_iw[0]~4_combout ;
wire \F_iw[0]~5_combout ;
wire \F_iw[0]~6_combout ;
wire \F_iw[0]~7_combout ;
wire \F_iw[0]~8_combout ;
wire \D_iw[0]~q ;
wire \F_iw[1]~9_combout ;
wire \F_iw[1]~10_combout ;
wire \F_iw[1]~11_combout ;
wire \F_iw[1]~12_combout ;
wire \D_iw[1]~q ;
wire \F_iw[4]~21_combout ;
wire \F_iw[4]~22_combout ;
wire \F_iw[4]~23_combout ;
wire \F_iw[4]~24_combout ;
wire \D_iw[4]~q ;
wire \F_iw[3]~17_combout ;
wire \F_iw[3]~18_combout ;
wire \F_iw[3]~19_combout ;
wire \F_iw[3]~20_combout ;
wire \D_iw[3]~q ;
wire \D_ctrl_ld_signed~0_combout ;
wire \D_ctrl_ld~2_combout ;
wire \D_ctrl_ld~3_combout ;
wire \R_ctrl_ld~q ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \Equal0~2_combout ;
wire \F_iw[5]~37_combout ;
wire \F_iw[5]~38_combout ;
wire \F_iw[5]~39_combout ;
wire \D_iw[5]~q ;
wire \Equal0~7_combout ;
wire \F_iw[15]~43_combout ;
wire \F_iw[15]~44_combout ;
wire \F_iw[15]~45_combout ;
wire \D_iw[15]~q ;
wire \D_ctrl_st~0_combout ;
wire \R_ctrl_st~q ;
wire \W_valid~3_combout ;
wire \W_valid~2_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \F_iw[14]~40_combout ;
wire \F_iw[14]~41_combout ;
wire \F_iw[14]~42_combout ;
wire \F_iw[14]~110_combout ;
wire \D_iw[14]~q ;
wire \D_op_opx_rsv63~0_combout ;
wire \F_iw[13]~28_combout ;
wire \F_iw[13]~29_combout ;
wire \F_iw[13]~30_combout ;
wire \D_iw[13]~q ;
wire \F_iw[16]~31_combout ;
wire \F_iw[16]~32_combout ;
wire \F_iw[16]~33_combout ;
wire \D_iw[16]~q ;
wire \F_iw[12]~34_combout ;
wire \F_iw[12]~35_combout ;
wire \F_iw[12]~36_combout ;
wire \D_iw[12]~q ;
wire \Equal62~4_combout ;
wire \Equal62~5_combout ;
wire \Equal62~6_combout ;
wire \D_ctrl_shift_rot~0_combout ;
wire \Equal62~7_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_shift_rot~3_combout ;
wire \R_ctrl_shift_rot~q ;
wire \E_shift_rot_cnt[0]~5_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~1_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \D_ctrl_alu_force_xor~14_combout ;
wire \Equal0~14_combout ;
wire \Equal0~15_combout ;
wire \D_dst_regnum[4]~3_combout ;
wire \Equal62~8_combout ;
wire \Equal62~14_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal62~12_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \Equal62~10_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \Equal0~13_combout ;
wire \Equal62~9_combout ;
wire \Equal0~3_combout ;
wire \D_op_cmpge~0_combout ;
wire \D_ctrl_exception~4_combout ;
wire \Equal62~11_combout ;
wire \D_op_opx_rsv17~0_combout ;
wire \D_ctrl_exception~5_combout ;
wire \Equal62~2_combout ;
wire \D_op_opx_rsv00~0_combout ;
wire \D_ctrl_exception~6_combout ;
wire \D_ctrl_exception~7_combout ;
wire \D_ctrl_exception~8_combout ;
wire \Equal0~11_combout ;
wire \D_ctrl_exception~9_combout ;
wire \D_ctrl_exception~10_combout ;
wire \Equal62~13_combout ;
wire \D_ctrl_exception~11_combout ;
wire \Equal62~3_combout ;
wire \Equal62~1_combout ;
wire \D_ctrl_exception~12_combout ;
wire \D_ctrl_exception~13_combout ;
wire \D_ctrl_exception~14_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \Equal0~4_combout ;
wire \Equal0~12_combout ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \D_ctrl_force_src2_zero~3_combout ;
wire \D_ctrl_force_src2_zero~4_combout ;
wire \D_ctrl_force_src2_zero~5_combout ;
wire \D_ctrl_force_src2_zero~6_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \R_src2_lo[4]~11_combout ;
wire \F_iw[6]~100_combout ;
wire \F_iw[6]~101_combout ;
wire \F_iw[6]~102_combout ;
wire \F_iw[6]~103_combout ;
wire \D_iw[6]~q ;
wire \D_dst_regnum[4]~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~5_combout ;
wire \Equal0~16_combout ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~1_combout ;
wire \D_ctrl_b_is_dst~2_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \R_ctrl_br_nxt~1_combout ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \E_src2[0]~16_combout ;
wire \R_src2_lo[0]~16_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~q ;
wire \E_shift_rot_cnt[0]~6 ;
wire \E_shift_rot_cnt[1]~7_combout ;
wire \F_iw[7]~96_combout ;
wire \F_iw[7]~97_combout ;
wire \F_iw[7]~98_combout ;
wire \F_iw[7]~99_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~15_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \E_shift_rot_cnt[1]~8 ;
wire \E_shift_rot_cnt[2]~9_combout ;
wire \F_iw[8]~89_combout ;
wire \F_iw[8]~90_combout ;
wire \F_iw[8]~91_combout ;
wire \F_iw[8]~92_combout ;
wire \D_iw[8]~q ;
wire \R_src2_lo[2]~14_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \E_shift_rot_cnt[2]~10 ;
wire \E_shift_rot_cnt[3]~11_combout ;
wire \F_iw[9]~83_combout ;
wire \F_iw[9]~84_combout ;
wire \F_iw[9]~85_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~13_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_shift_rot_cnt[3]~12 ;
wire \E_shift_rot_cnt[4]~13_combout ;
wire \F_iw[10]~77_combout ;
wire \F_iw[10]~78_combout ;
wire \F_iw[10]~79_combout ;
wire \D_iw[10]~q ;
wire \R_src2_lo[4]~12_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~0_combout ;
wire \E_stall~1_combout ;
wire \E_stall~2_combout ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data~q ;
wire \D_ctrl_mem16~0_combout ;
wire \av_ld_align_cycle_nxt[0]~0_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \av_ld_align_cycle_nxt[1]~1_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \av_ld_aligning_data_nxt~2_combout ;
wire \E_stall~3_combout ;
wire \E_stall~4_combout ;
wire \E_valid_from_R~3_combout ;
wire \E_valid_from_R~2_combout ;
wire \E_valid_from_R~q ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \D_ctrl_jmp_direct~1_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_ctrl_br~q ;
wire \D_ctrl_retaddr~4_combout ;
wire \D_ctrl_retaddr~5_combout ;
wire \D_ctrl_retaddr~6_combout ;
wire \Equal0~9_combout ;
wire \D_ctrl_retaddr~7_combout ;
wire \D_ctrl_retaddr~8_combout ;
wire \D_ctrl_retaddr~9_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~11_combout ;
wire \R_src1[1]~12_combout ;
wire \E_src1[1]~q ;
wire \D_op_wrctl~combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \W_ienable_reg_nxt~0_combout ;
wire \W_ienable_reg_nxt~1_combout ;
wire \W_ienable_reg[1]~q ;
wire \W_ipending_reg_nxt[1]~0_combout ;
wire \W_ipending_reg[1]~q ;
wire \R_src1[0]~13_combout ;
wire \E_src1[0]~q ;
wire \W_ienable_reg[0]~q ;
wire \W_ipending_reg_nxt[0]~1_combout ;
wire \W_ipending_reg[0]~q ;
wire \D_ctrl_exception~0_combout ;
wire \D_ctrl_exception~1_combout ;
wire \D_ctrl_exception~2_combout ;
wire \D_ctrl_exception~3_combout ;
wire \D_dst_regnum[4]~1_combout ;
wire \D_dst_regnum[4]~2_combout ;
wire \D_dst_regnum[4]~4_combout ;
wire \D_ctrl_exception~15_combout ;
wire \R_ctrl_exception~q ;
wire \D_ctrl_break~0_combout ;
wire \R_ctrl_break~q ;
wire \F_pc_no_crst_nxt[25]~5_combout ;
wire \Equal132~2_combout ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \W_estatus_reg_inst_nxt~1_combout ;
wire \W_estatus_reg~q ;
wire \Equal132~1_combout ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \W_bstatus_reg_inst_nxt~1_combout ;
wire \W_bstatus_reg~q ;
wire \Equal132~0_combout ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \D_op_eret~combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_status_reg_pie~q ;
wire \D_iw[26]~0_combout ;
wire \D_iw[26]~1_combout ;
wire \F_iw[11]~25_combout ;
wire \F_iw[11]~26_combout ;
wire \F_iw[11]~27_combout ;
wire \D_iw[11]~q ;
wire \Equal62~0_combout ;
wire \Equal0~5_combout ;
wire \D_ctrl_alu_subtract~8_combout ;
wire \D_ctrl_alu_subtract~9_combout ;
wire \D_ctrl_alu_subtract~5_combout ;
wire \D_ctrl_alu_subtract~10_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \F_iw[21]~46_combout ;
wire \F_iw[21]~47_combout ;
wire \F_iw[21]~48_combout ;
wire \D_iw[21]~q ;
wire \E_src2[28]~0_combout ;
wire \F_iw[18]~49_combout ;
wire \F_iw[18]~50_combout ;
wire \F_iw[18]~51_combout ;
wire \F_iw[18]~52_combout ;
wire \D_iw[18]~q ;
wire \Equal0~6_combout ;
wire \D_ctrl_unsigned_lo_imm16~3_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~4_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi~0_combout ;
wire \E_src2[28]~q ;
wire \Add1~0_combout ;
wire \R_src1~10_combout ;
wire \E_src1[28]~0_combout ;
wire \F_pc_plus_one[0]~1 ;
wire \F_pc_plus_one[1]~3 ;
wire \F_pc_plus_one[2]~5 ;
wire \F_pc_plus_one[3]~7 ;
wire \F_pc_plus_one[4]~9 ;
wire \F_pc_plus_one[5]~11 ;
wire \F_pc_plus_one[6]~13 ;
wire \F_pc_plus_one[7]~15 ;
wire \F_pc_plus_one[8]~17 ;
wire \F_pc_plus_one[9]~19 ;
wire \F_pc_plus_one[10]~21 ;
wire \F_pc_plus_one[11]~23 ;
wire \F_pc_plus_one[12]~25 ;
wire \F_pc_plus_one[13]~27 ;
wire \F_pc_plus_one[14]~29 ;
wire \F_pc_plus_one[15]~31 ;
wire \F_pc_plus_one[16]~33 ;
wire \F_pc_plus_one[17]~35 ;
wire \F_pc_plus_one[18]~37 ;
wire \F_pc_plus_one[19]~39 ;
wire \F_pc_plus_one[20]~41 ;
wire \F_pc_plus_one[21]~43 ;
wire \F_pc_plus_one[22]~45 ;
wire \F_pc_plus_one[23]~47 ;
wire \F_pc_plus_one[24]~49 ;
wire \F_pc_plus_one[25]~51 ;
wire \F_pc_plus_one[26]~52_combout ;
wire \E_src1[28]~q ;
wire \E_src2[27]~1_combout ;
wire \F_iw[17]~53_combout ;
wire \F_iw[17]~54_combout ;
wire \F_iw[17]~55_combout ;
wire \F_iw[17]~111_combout ;
wire \D_iw[17]~q ;
wire \E_src2[27]~q ;
wire \Add1~1_combout ;
wire \F_iw[31]~56_combout ;
wire \F_iw[31]~57_combout ;
wire \F_iw[31]~58_combout ;
wire \D_iw[31]~q ;
wire \E_src1[27]~1_combout ;
wire \F_pc_plus_one[25]~50_combout ;
wire \E_src1[27]~q ;
wire \E_src2[26]~2_combout ;
wire \E_src2[26]~q ;
wire \Add1~2_combout ;
wire \F_iw[30]~59_combout ;
wire \F_iw[30]~60_combout ;
wire \F_iw[30]~61_combout ;
wire \D_iw[30]~q ;
wire \E_src1[26]~2_combout ;
wire \F_pc_plus_one[24]~48_combout ;
wire \E_src1[26]~q ;
wire \E_src2[25]~3_combout ;
wire \E_src2[25]~q ;
wire \Add1~3_combout ;
wire \F_iw[29]~62_combout ;
wire \F_iw[29]~63_combout ;
wire \F_iw[29]~64_combout ;
wire \D_iw[29]~q ;
wire \E_src1[25]~3_combout ;
wire \F_pc_plus_one[23]~46_combout ;
wire \E_src1[25]~q ;
wire \E_src2[24]~4_combout ;
wire \E_src2[24]~q ;
wire \Add1~4_combout ;
wire \F_iw[28]~65_combout ;
wire \F_iw[28]~66_combout ;
wire \F_iw[28]~67_combout ;
wire \D_iw[28]~q ;
wire \E_src1[24]~4_combout ;
wire \F_pc_plus_one[22]~44_combout ;
wire \E_src1[24]~q ;
wire \E_src2[23]~5_combout ;
wire \E_src2[23]~q ;
wire \Add1~5_combout ;
wire \F_iw[27]~68_combout ;
wire \F_iw[27]~69_combout ;
wire \F_iw[27]~70_combout ;
wire \D_iw[27]~q ;
wire \E_src1[23]~5_combout ;
wire \F_pc_plus_one[21]~42_combout ;
wire \E_src1[23]~q ;
wire \E_src2[22]~6_combout ;
wire \E_src2[22]~q ;
wire \Add1~6_combout ;
wire \F_iw[26]~71_combout ;
wire \F_iw[26]~72_combout ;
wire \F_iw[26]~73_combout ;
wire \D_iw[26]~q ;
wire \E_src1[22]~6_combout ;
wire \F_pc_plus_one[20]~40_combout ;
wire \E_src1[22]~q ;
wire \E_src2[21]~7_combout ;
wire \E_src2[21]~q ;
wire \Add1~7_combout ;
wire \F_iw[25]~74_combout ;
wire \F_iw[25]~75_combout ;
wire \F_iw[25]~76_combout ;
wire \D_iw[25]~q ;
wire \E_src1[21]~7_combout ;
wire \F_pc_plus_one[19]~38_combout ;
wire \E_src1[21]~q ;
wire \E_src2[20]~8_combout ;
wire \E_src2[20]~q ;
wire \Add1~8_combout ;
wire \F_iw[24]~80_combout ;
wire \F_iw[24]~81_combout ;
wire \F_iw[24]~82_combout ;
wire \D_iw[24]~q ;
wire \E_src1[20]~8_combout ;
wire \F_pc_plus_one[18]~36_combout ;
wire \E_src1[20]~q ;
wire \E_src2[19]~9_combout ;
wire \E_src2[19]~q ;
wire \Add1~9_combout ;
wire \F_iw[23]~86_combout ;
wire \F_iw[23]~87_combout ;
wire \F_iw[23]~88_combout ;
wire \D_iw[23]~q ;
wire \E_src1[19]~9_combout ;
wire \F_pc_plus_one[17]~34_combout ;
wire \E_src1[19]~q ;
wire \E_src2[18]~10_combout ;
wire \E_src2[18]~q ;
wire \Add1~10_combout ;
wire \F_iw[22]~93_combout ;
wire \F_iw[22]~94_combout ;
wire \F_iw[22]~95_combout ;
wire \D_iw[22]~q ;
wire \E_src1[18]~10_combout ;
wire \F_pc_plus_one[16]~32_combout ;
wire \E_src1[18]~q ;
wire \E_src2[17]~11_combout ;
wire \E_src2[17]~q ;
wire \Add1~11_combout ;
wire \E_src1[17]~11_combout ;
wire \F_pc_plus_one[15]~30_combout ;
wire \E_src1[17]~q ;
wire \E_src2[16]~12_combout ;
wire \E_src2[16]~q ;
wire \Add1~12_combout ;
wire \F_iw[20]~104_combout ;
wire \F_iw[20]~105_combout ;
wire \F_iw[20]~106_combout ;
wire \D_iw[20]~q ;
wire \E_src1[16]~12_combout ;
wire \F_pc_plus_one[14]~28_combout ;
wire \E_src1[16]~q ;
wire \E_src2[5]~15_combout ;
wire \R_src2_lo[15]~0_combout ;
wire \E_src2[15]~q ;
wire \Add1~13_combout ;
wire \F_iw[19]~107_combout ;
wire \F_iw[19]~108_combout ;
wire \F_iw[19]~109_combout ;
wire \D_iw[19]~q ;
wire \E_src1[15]~13_combout ;
wire \F_pc_plus_one[13]~26_combout ;
wire \E_src1[15]~q ;
wire \R_src2_lo[14]~1_combout ;
wire \E_src2[14]~q ;
wire \Add1~14_combout ;
wire \E_src1[14]~14_combout ;
wire \F_pc_plus_one[12]~24_combout ;
wire \E_src1[14]~q ;
wire \R_src2_lo[13]~2_combout ;
wire \E_src2[13]~q ;
wire \Add1~15_combout ;
wire \E_src1[13]~15_combout ;
wire \F_pc_plus_one[11]~22_combout ;
wire \E_src1[13]~q ;
wire \R_src2_lo[12]~3_combout ;
wire \E_src2[12]~q ;
wire \Add1~16_combout ;
wire \E_src1[12]~16_combout ;
wire \F_pc_plus_one[10]~20_combout ;
wire \E_src1[12]~q ;
wire \R_src2_lo[11]~4_combout ;
wire \E_src2[11]~q ;
wire \Add1~17_combout ;
wire \E_src1[11]~17_combout ;
wire \F_pc_plus_one[9]~18_combout ;
wire \E_src1[11]~q ;
wire \R_src2_lo[10]~5_combout ;
wire \E_src2[10]~q ;
wire \Add1~18_combout ;
wire \E_src1[10]~18_combout ;
wire \F_pc_plus_one[8]~16_combout ;
wire \E_src1[10]~q ;
wire \R_src2_lo[9]~6_combout ;
wire \E_src2[9]~q ;
wire \Add1~19_combout ;
wire \E_src1[9]~19_combout ;
wire \F_pc_plus_one[7]~14_combout ;
wire \E_src1[9]~q ;
wire \R_src2_lo[8]~7_combout ;
wire \E_src2[8]~q ;
wire \Add1~20_combout ;
wire \E_src1[8]~20_combout ;
wire \F_pc_plus_one[6]~12_combout ;
wire \E_src1[8]~q ;
wire \R_src2_lo[7]~8_combout ;
wire \E_src2[7]~q ;
wire \Add1~21_combout ;
wire \E_src1[7]~21_combout ;
wire \F_pc_plus_one[5]~10_combout ;
wire \E_src1[7]~q ;
wire \R_src2_lo[6]~9_combout ;
wire \E_src2[6]~q ;
wire \Add1~22_combout ;
wire \E_src1[6]~22_combout ;
wire \F_pc_plus_one[4]~8_combout ;
wire \E_src1[6]~q ;
wire \R_src2_lo[5]~10_combout ;
wire \E_src2[5]~q ;
wire \Add1~23_combout ;
wire \E_src1[5]~23_combout ;
wire \F_pc_plus_one[3]~6_combout ;
wire \E_src1[5]~q ;
wire \Add1~24_combout ;
wire \E_src1[4]~24_combout ;
wire \F_pc_plus_one[2]~4_combout ;
wire \E_src1[4]~q ;
wire \Add1~25_combout ;
wire \E_src1[3]~26_combout ;
wire \F_pc_plus_one[1]~2_combout ;
wire \E_src1[3]~q ;
wire \Add1~26_combout ;
wire \E_src1[2]~25_combout ;
wire \F_pc_plus_one[0]~0_combout ;
wire \E_src1[2]~q ;
wire \Add1~27_combout ;
wire \Add1~28_combout ;
wire \Add1~30_cout ;
wire \Add1~32 ;
wire \Add1~34 ;
wire \Add1~36 ;
wire \Add1~38 ;
wire \Add1~40 ;
wire \Add1~42 ;
wire \Add1~44 ;
wire \Add1~46 ;
wire \Add1~48 ;
wire \Add1~50 ;
wire \Add1~52 ;
wire \Add1~54 ;
wire \Add1~56 ;
wire \Add1~58 ;
wire \Add1~60 ;
wire \Add1~62 ;
wire \Add1~64 ;
wire \Add1~66 ;
wire \Add1~68 ;
wire \Add1~70 ;
wire \Add1~72 ;
wire \Add1~74 ;
wire \Add1~76 ;
wire \Add1~78 ;
wire \Add1~80 ;
wire \Add1~82 ;
wire \Add1~84 ;
wire \Add1~86 ;
wire \Add1~87_combout ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~10_combout ;
wire \D_ctrl_alu_force_xor~11_combout ;
wire \D_ctrl_alu_force_xor~13_combout ;
wire \D_ctrl_alu_force_xor~12_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[28]~0_combout ;
wire \Equal0~8_combout ;
wire \D_ctrl_logic~combout ;
wire \R_ctrl_logic~q ;
wire \W_alu_result[28]~0_combout ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \E_shift_rot_result_nxt[27]~1_combout ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[26]~2_combout ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[25]~3_combout ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[24]~4_combout ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[23]~5_combout ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[22]~6_combout ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[21]~7_combout ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[20]~8_combout ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[19]~9_combout ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[18]~10_combout ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[17]~11_combout ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[16]~12_combout ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[15]~13_combout ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[14]~14_combout ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[13]~15_combout ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[12]~20_combout ;
wire \E_shift_rot_result[12]~q ;
wire \E_shift_rot_result_nxt[11]~24_combout ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[10]~21_combout ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[9]~22_combout ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[8]~23_combout ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[7]~17_combout ;
wire \E_shift_rot_result[7]~q ;
wire \E_shift_rot_result_nxt[6]~16_combout ;
wire \E_shift_rot_result[6]~q ;
wire \E_shift_rot_result_nxt[5]~18_combout ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[4]~19_combout ;
wire \E_shift_rot_result[4]~q ;
wire \E_shift_rot_result_nxt[3]~26_combout ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[2]~25_combout ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[1]~28_combout ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[0]~30_combout ;
wire \E_shift_rot_result[0]~q ;
wire \R_ctrl_rot_right_nxt~0_combout ;
wire \R_ctrl_rot_right~q ;
wire \D_ctrl_shift_logical~1_combout ;
wire \D_ctrl_shift_logical~2_combout ;
wire \R_ctrl_shift_logical~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[31]~31_combout ;
wire \R_src1[31]~14_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_result_nxt[30]~29_combout ;
wire \R_src1[30]~15_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[29]~27_combout ;
wire \R_src1[29]~16_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[28]~0_combout ;
wire \E_shift_rot_result[28]~q ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \D_ctrl_br_cmp~2_combout ;
wire \D_ctrl_br_cmp~5_combout ;
wire \D_ctrl_br_cmp~3_combout ;
wire \D_ctrl_br_cmp~4_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~0_combout ;
wire \Add1~85_combout ;
wire \E_logic_result[27]~1_combout ;
wire \W_alu_result[27]~1_combout ;
wire \Add1~83_combout ;
wire \E_logic_result[26]~2_combout ;
wire \W_alu_result[26]~2_combout ;
wire \Add1~81_combout ;
wire \E_logic_result[25]~3_combout ;
wire \W_alu_result[25]~3_combout ;
wire \Add1~79_combout ;
wire \E_logic_result[24]~4_combout ;
wire \W_alu_result[24]~4_combout ;
wire \Add1~77_combout ;
wire \E_logic_result[23]~5_combout ;
wire \W_alu_result[23]~5_combout ;
wire \Add1~75_combout ;
wire \E_logic_result[22]~6_combout ;
wire \W_alu_result[22]~6_combout ;
wire \Add1~73_combout ;
wire \E_logic_result[21]~7_combout ;
wire \W_alu_result[21]~7_combout ;
wire \Add1~71_combout ;
wire \E_logic_result[20]~8_combout ;
wire \W_alu_result[20]~8_combout ;
wire \Add1~69_combout ;
wire \E_logic_result[19]~9_combout ;
wire \W_alu_result[19]~9_combout ;
wire \Add1~67_combout ;
wire \E_logic_result[18]~10_combout ;
wire \W_alu_result[18]~10_combout ;
wire \Add1~65_combout ;
wire \E_logic_result[17]~11_combout ;
wire \W_alu_result[17]~11_combout ;
wire \Add1~63_combout ;
wire \E_logic_result[16]~12_combout ;
wire \W_alu_result[16]~12_combout ;
wire \Add1~61_combout ;
wire \E_logic_result[15]~13_combout ;
wire \W_alu_result[15]~13_combout ;
wire \Add1~59_combout ;
wire \E_logic_result[14]~14_combout ;
wire \W_alu_result[14]~14_combout ;
wire \Add1~57_combout ;
wire \E_logic_result[13]~15_combout ;
wire \W_alu_result[13]~15_combout ;
wire \Add1~43_combout ;
wire \E_logic_result[6]~16_combout ;
wire \W_alu_result[6]~22_combout ;
wire \Add1~45_combout ;
wire \E_logic_result[7]~17_combout ;
wire \W_alu_result[7]~21_combout ;
wire \Add1~41_combout ;
wire \E_logic_result[5]~18_combout ;
wire \W_alu_result[5]~23_combout ;
wire \Add1~39_combout ;
wire \E_logic_result[4]~19_combout ;
wire \W_alu_result[4]~24_combout ;
wire \Add1~55_combout ;
wire \E_logic_result[12]~20_combout ;
wire \W_alu_result[12]~16_combout ;
wire \Add1~51_combout ;
wire \E_logic_result[10]~21_combout ;
wire \W_alu_result[10]~18_combout ;
wire \Add1~49_combout ;
wire \E_logic_result[9]~22_combout ;
wire \W_alu_result[9]~19_combout ;
wire \Add1~47_combout ;
wire \E_logic_result[8]~23_combout ;
wire \W_alu_result[8]~20_combout ;
wire \Add1~53_combout ;
wire \E_logic_result[11]~24_combout ;
wire \W_alu_result[11]~17_combout ;
wire \Add1~35_combout ;
wire \E_logic_result[2]~25_combout ;
wire \W_alu_result[2]~25_combout ;
wire \Add1~37_combout ;
wire \E_logic_result[3]~26_combout ;
wire \W_alu_result[3]~26_combout ;
wire \D_ctrl_mem16~1_combout ;
wire \d_writedata[31]~3_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \d_writedata[30]~4_combout ;
wire \d_writedata[29]~5_combout ;
wire \d_writedata[28]~6_combout ;
wire \d_writedata[27]~7_combout ;
wire \d_writedata[26]~2_combout ;
wire \d_writedata[25]~1_combout ;
wire \d_writedata[24]~0_combout ;
wire \d_read_nxt~0_combout ;
wire \E_st_stall~combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_uncond_cti_non_br~2_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~19_combout ;
wire \R_ctrl_br_uncond~q ;
wire \R_compare_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \R_compare_op[0]~q ;
wire \Equal127~0_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \Equal127~3_combout ;
wire \Equal127~4_combout ;
wire \Equal127~5_combout ;
wire \Equal127~6_combout ;
wire \R_src2_hi[15]~1_combout ;
wire \R_src2_hi[15]~2_combout ;
wire \E_src2[31]~q ;
wire \E_logic_result[31]~27_combout ;
wire \Equal127~7_combout ;
wire \E_src2[30]~13_combout ;
wire \E_src2[30]~q ;
wire \E_logic_result[30]~28_combout ;
wire \E_src2[29]~14_combout ;
wire \E_src2[29]~q ;
wire \E_logic_result[29]~29_combout ;
wire \E_logic_result[1]~30_combout ;
wire \E_logic_result[0]~31_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \E_cmp_result~0_combout ;
wire \E_invert_arith_src_msb~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~q ;
wire \Add1~89_combout ;
wire \E_arith_src1[31]~combout ;
wire \Add1~90_combout ;
wire \Add1~91_combout ;
wire \Add1~88 ;
wire \Add1~93 ;
wire \Add1~95 ;
wire \Add1~97 ;
wire \Add1~98_combout ;
wire \E_cmp_result~1_combout ;
wire \W_cmp_result~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_no_crst_nxt[26]~32_combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \F_pc_no_crst_nxt[26]~4_combout ;
wire \F_pc_no_crst_nxt[25]~6_combout ;
wire \F_pc_no_crst_nxt[24]~7_combout ;
wire \F_pc_no_crst_nxt[23]~8_combout ;
wire \F_pc_no_crst_nxt[22]~9_combout ;
wire \F_pc_no_crst_nxt[21]~10_combout ;
wire \F_pc_no_crst_nxt[20]~11_combout ;
wire \F_pc_no_crst_nxt[19]~12_combout ;
wire \F_pc_no_crst_nxt[18]~13_combout ;
wire \F_pc_no_crst_nxt[17]~14_combout ;
wire \F_pc_no_crst_nxt[16]~15_combout ;
wire \F_pc_no_crst_nxt[15]~16_combout ;
wire \F_pc_no_crst_nxt[14]~17_combout ;
wire \F_pc_no_crst_nxt[13]~18_combout ;
wire \F_pc_no_crst_nxt[12]~19_combout ;
wire \F_pc_no_crst_nxt[11]~20_combout ;
wire \F_pc_no_crst_nxt[10]~33_combout ;
wire \F_pc_no_crst_nxt[10]~21_combout ;
wire \F_pc_no_crst_nxt[8]~22_combout ;
wire \F_pc_no_crst_nxt[7]~23_combout ;
wire \F_pc_no_crst_nxt[6]~24_combout ;
wire \F_pc_no_crst_nxt[5]~25_combout ;
wire \F_pc_no_crst_nxt[3]~26_combout ;
wire \i_read_nxt~0_combout ;
wire \F_pc_no_crst_nxt[2]~27_combout ;
wire \F_pc_no_crst_nxt[4]~28_combout ;
wire \F_pc_no_crst_nxt[9]~29_combout ;
wire \Add1~31_combout ;
wire \Add1~33_combout ;
wire \E_mem_byte_en[0]~0_combout ;
wire \F_pc_no_crst_nxt[0]~30_combout ;
wire \F_pc_no_crst_nxt[1]~31_combout ;
wire \E_st_data[8]~0_combout ;
wire \E_st_data[9]~1_combout ;
wire \E_st_data[10]~2_combout ;
wire \E_st_data[11]~3_combout ;
wire \E_st_data[12]~4_combout ;
wire \E_st_data[13]~5_combout ;
wire \E_st_data[14]~6_combout ;
wire \E_st_data[15]~7_combout ;
wire \d_writedata[22]~8_combout ;
wire \E_st_data[16]~8_combout ;
wire \E_st_data[17]~9_combout ;
wire \hbreak_enabled~0_combout ;
wire \E_mem_byte_en[2]~1_combout ;
wire \E_mem_byte_en[1]~2_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \E_st_data[21]~10_combout ;
wire \E_st_data[18]~11_combout ;
wire \E_st_data[23]~12_combout ;
wire \E_st_data[22]~13_combout ;
wire \E_st_data[20]~14_combout ;
wire \E_st_data[19]~15_combout ;


final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_oci the_final_project_soc_nios2_qsys_0_cpu_nios2_oci(
	.sr_0(sr_0),
	.jtag_break(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|jtag_break~q ),
	.readdata_0(readdata_01),
	.readdata_1(readdata_11),
	.readdata_2(readdata_21),
	.readdata_3(readdata_3),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr1(WideOr11),
	.local_read(local_read),
	.hbreak_enabled(hbreak_enabled1),
	.mem(mem),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_411,src_data_40,src_data_39,src_data_38}),
	.oci_ienable_1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.oci_ienable_0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_single_step_mode(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.r_early_rst(r_early_rst),
	.readdata_4(readdata_41),
	.readdata_11(readdata_111),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_5(readdata_5),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_21(readdata_211),
	.readdata_18(readdata_18),
	.readdata_17(readdata_171),
	.readdata_31(readdata_311),
	.readdata_30(readdata_30),
	.readdata_29(readdata_29),
	.readdata_28(readdata_28),
	.readdata_27(readdata_27),
	.readdata_26(readdata_26),
	.readdata_25(readdata_25),
	.readdata_10(readdata_10),
	.readdata_24(readdata_24),
	.readdata_9(readdata_9),
	.readdata_23(readdata_23),
	.readdata_8(readdata_81),
	.readdata_22(readdata_22),
	.readdata_7(readdata_71),
	.readdata_6(readdata_61),
	.readdata_20(readdata_20),
	.readdata_19(readdata_19),
	.debugaccess_nxt(src_payload7),
	.writedata_nxt({src_payload23,src_payload24,src_payload25,src_payload26,src_payload27,src_payload28,src_payload29,src_payload31,src_payload33,src_payload35,src_payload20,src_payload38,src_payload39,src_payload21,src_payload22,src_payload15,src_payload19,src_payload18,src_payload14,
src_payload16,src_payload13,src_payload30,src_payload32,src_payload34,src_payload36,src_payload37,src_payload17,src_payload12,src_payload10,src_payload11,src_payload9,src_payload8}),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_register_bank_b_module final_project_soc_nios2_qsys_0_cpu_register_bank_b(
	.q_b_0(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_8(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_9(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_10(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_11(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_12(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_15(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_16(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_17(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_28(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_31(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.D_iw_26(\D_iw[26]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_22(\D_iw[22]~q ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~4_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~5_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~6_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~7_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~8_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~9_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~10_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~11_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~12_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~13_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~14_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~15_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~16_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~17_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~18_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~19_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~20_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~21_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~22_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~23_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~24_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~25_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~26_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~27_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~28_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~29_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~30_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~31_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~32_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~33_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~34_combout ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_register_bank_a_module final_project_soc_nios2_qsys_0_cpu_register_bank_a(
	.q_b_28(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_1(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_31(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.D_iw_31(\D_iw[31]~q ),
	.D_iw_30(\D_iw[30]~q ),
	.D_iw_29(\D_iw[29]~q ),
	.D_iw_28(\D_iw[28]~q ),
	.D_iw_27(\D_iw[27]~q ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~4_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~5_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~6_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~7_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~8_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~9_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~10_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~11_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~12_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~13_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~14_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~15_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~16_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~17_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~18_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~19_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~20_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~21_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~22_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~23_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~24_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~25_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~26_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~27_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~28_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~29_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~30_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~31_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~32_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~33_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~34_combout ),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \Add1~92 (
	.dataa(\Add1~91_combout ),
	.datab(\E_src1[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~88 ),
	.combout(\Add1~92_combout ),
	.cout(\Add1~93 ));
defparam \Add1~92 .lut_mask = 16'h96EF;
defparam \Add1~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~94 (
	.dataa(\Add1~90_combout ),
	.datab(\E_src1[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~93 ),
	.combout(\Add1~94_combout ),
	.cout(\Add1~95 ));
defparam \Add1~94 .lut_mask = 16'h967F;
defparam \Add1~94 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~96 (
	.dataa(\Add1~89_combout ),
	.datab(\E_arith_src1[31]~combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~95 ),
	.combout(\Add1~96_combout ),
	.cout(\Add1~97 ));
defparam \Add1~96 .lut_mask = 16'h96EF;
defparam \Add1~96 .sum_lutc_input = "cin";

dffeas \W_alu_result[0] (
	.clk(clk_clk),
	.d(\W_alu_result[0]~27_combout ),
	.asdata(\E_shift_rot_result[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

dffeas \W_alu_result[1] (
	.clk(clk_clk),
	.d(\W_alu_result[1]~28_combout ),
	.asdata(\E_shift_rot_result[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

dffeas \av_ld_byte1_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[0]~0_combout ),
	.asdata(\av_ld_byte2_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

dffeas \av_ld_byte1_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[1]~1_combout ),
	.asdata(\av_ld_byte2_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

dffeas \av_ld_byte1_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[2]~2_combout ),
	.asdata(\av_ld_byte2_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

dffeas \av_ld_byte1_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[3]~3_combout ),
	.asdata(\av_ld_byte2_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

dffeas \av_ld_byte1_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[4]~4_combout ),
	.asdata(\av_ld_byte2_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

dffeas \av_ld_byte1_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[5]~5_combout ),
	.asdata(\av_ld_byte2_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

dffeas \av_ld_byte1_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[6]~6_combout ),
	.asdata(\av_ld_byte2_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

dffeas \av_ld_byte1_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[7]~7_combout ),
	.asdata(\av_ld_byte2_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

dffeas \av_ld_byte2_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[0]~0_combout ),
	.asdata(\av_ld_byte3_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

dffeas \av_ld_byte2_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[1]~1_combout ),
	.asdata(\av_ld_byte3_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

dffeas \av_ld_byte2_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[7]~2_combout ),
	.asdata(\av_ld_byte3_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

dffeas \av_ld_byte2_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[6]~3_combout ),
	.asdata(\av_ld_byte3_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

dffeas \av_ld_byte2_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[5]~4_combout ),
	.asdata(\av_ld_byte3_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

dffeas \av_ld_byte2_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[4]~5_combout ),
	.asdata(\av_ld_byte3_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

dffeas \av_ld_byte2_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[3]~6_combout ),
	.asdata(\av_ld_byte3_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

dffeas \av_ld_byte2_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[2]~7_combout ),
	.asdata(\av_ld_byte3_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

cycloneive_lcell_comb \W_alu_result[0]~27 (
	.dataa(\Add1~31_combout ),
	.datab(\E_logic_result[0]~31_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[0]~27_combout ),
	.cout());
defparam \W_alu_result[0]~27 .lut_mask = 16'hAACC;
defparam \W_alu_result[0]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[1]~28 (
	.dataa(\Add1~33_combout ),
	.datab(\E_logic_result[1]~30_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[1]~28_combout ),
	.cout());
defparam \W_alu_result[1]~28 .lut_mask = 16'hAACC;
defparam \W_alu_result[1]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[0]~0 (
	.dataa(src_data_8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte1_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[1]~1 (
	.dataa(src_data_9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[1]~1_combout ),
	.cout());
defparam \av_ld_byte1_data[1]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[2]~2 (
	.dataa(src_data_10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[2]~2_combout ),
	.cout());
defparam \av_ld_byte1_data[2]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[3]~3 (
	.dataa(src_data_111),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[3]~3_combout ),
	.cout());
defparam \av_ld_byte1_data[3]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[4]~4 (
	.dataa(src_data_12),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[4]~4_combout ),
	.cout());
defparam \av_ld_byte1_data[4]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[5]~5 (
	.dataa(src_data_13),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[5]~5_combout ),
	.cout());
defparam \av_ld_byte1_data[5]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[6]~6 (
	.dataa(src_data_14),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[6]~6_combout ),
	.cout());
defparam \av_ld_byte1_data[6]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[7]~7 (
	.dataa(src_data_15),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[7]~7_combout ),
	.cout());
defparam \av_ld_byte1_data[7]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[0]~0 (
	.dataa(src_data_16),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte2_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[1]~1 (
	.dataa(src_data_17),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[1]~1_combout ),
	.cout());
defparam \av_ld_byte2_data[1]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[7]~2 (
	.dataa(src_data_23),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[7]~2_combout ),
	.cout());
defparam \av_ld_byte2_data[7]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[7]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[6]~3 (
	.dataa(src_data_22),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[6]~3_combout ),
	.cout());
defparam \av_ld_byte2_data[6]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[6]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[5]~4 (
	.dataa(src_data_211),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[5]~4_combout ),
	.cout());
defparam \av_ld_byte2_data[5]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[5]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[4]~5 (
	.dataa(src_data_20),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[4]~5_combout ),
	.cout());
defparam \av_ld_byte2_data[4]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[3]~6 (
	.dataa(src_data_19),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[3]~6_combout ),
	.cout());
defparam \av_ld_byte2_data[3]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[3]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[2]~7 (
	.dataa(src_data_18),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[2]~7_combout ),
	.cout());
defparam \av_ld_byte2_data[2]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[2]~7 .sum_lutc_input = "datac";

dffeas \W_alu_result[31] (
	.clk(clk_clk),
	.d(\W_alu_result[31]~29_combout ),
	.asdata(\E_shift_rot_result[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(clk_clk),
	.d(\W_alu_result[30]~30_combout ),
	.asdata(\E_shift_rot_result[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(clk_clk),
	.d(\W_alu_result[29]~31_combout ),
	.asdata(\E_shift_rot_result[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

cycloneive_lcell_comb \W_alu_result[31]~29 (
	.dataa(\Add1~96_combout ),
	.datab(\E_logic_result[31]~27_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[31]~29_combout ),
	.cout());
defparam \W_alu_result[31]~29 .lut_mask = 16'hAACC;
defparam \W_alu_result[31]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[30]~30 (
	.dataa(\Add1~94_combout ),
	.datab(\E_logic_result[30]~28_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[30]~30_combout ),
	.cout());
defparam \W_alu_result[30]~30 .lut_mask = 16'hAACC;
defparam \W_alu_result[30]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[29]~31 (
	.dataa(\Add1~92_combout ),
	.datab(\E_logic_result[29]~29_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[29]~31_combout ),
	.cout());
defparam \W_alu_result[29]~31 .lut_mask = 16'hAACC;
defparam \W_alu_result[29]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld_signed~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~1_combout ),
	.cout());
defparam \D_ctrl_ld_signed~1 .lut_mask = 16'hEEEE;
defparam \D_ctrl_ld_signed~1 .sum_lutc_input = "datac";

dffeas R_wr_dst_reg(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cycloneive_lcell_comb W_rf_wren(
	.dataa(r_sync_rst),
	.datab(\W_valid~q ),
	.datac(\R_wr_dst_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wren~combout ),
	.cout());
defparam W_rf_wren.lut_mask = 16'hFEFE;
defparam W_rf_wren.sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[0]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~0 (
	.dataa(\W_cmp_result~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~0_combout ),
	.cout());
defparam \W_rf_wr_data[0]~0 .lut_mask = 16'hEEEE;
defparam \W_rf_wr_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_control_rd_data[0] (
	.clk(clk_clk),
	.d(\E_control_rd_data[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~1 (
	.dataa(\W_control_rd_data[0]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~1_combout ),
	.cout());
defparam \W_rf_wr_data[0]~1 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[0]~2 (
	.dataa(\av_ld_byte0_data[0]~q ),
	.datab(\W_rf_wr_data[0]~0_combout ),
	.datac(\W_rf_wr_data[0]~1_combout ),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~2_combout ),
	.cout());
defparam \W_rf_wr_data[0]~2 .lut_mask = 16'hFAFC;
defparam \W_rf_wr_data[0]~2 .sum_lutc_input = "datac";

dffeas \R_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

dffeas \av_ld_byte0_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

dffeas \W_control_rd_data[1] (
	.clk(clk_clk),
	.d(\E_control_rd_data[1]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[1]~q ),
	.prn(vcc));
defparam \W_control_rd_data[1] .is_wysiwyg = "true";
defparam \W_control_rd_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[1]~3 (
	.dataa(\W_control_rd_data[1]~q ),
	.datab(\W_alu_result[1]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~3_combout ),
	.cout());
defparam \W_rf_wr_data[1]~3 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[1]~4 (
	.dataa(\av_ld_byte0_data[1]~q ),
	.datab(\W_rf_wr_data[1]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~4_combout ),
	.cout());
defparam \W_rf_wr_data[1]~4 .lut_mask = 16'hAACC;
defparam \W_rf_wr_data[1]~4 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[2]~5 (
	.dataa(\av_ld_byte0_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_2),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[2]~5_combout ),
	.cout());
defparam \W_rf_wr_data[2]~5 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[2]~5 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[3]~6 (
	.dataa(\av_ld_byte0_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_3),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[3]~6_combout ),
	.cout());
defparam \W_rf_wr_data[3]~6 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[3]~6 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[4]~7 (
	.dataa(\av_ld_byte0_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_4),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[4]~7_combout ),
	.cout());
defparam \W_rf_wr_data[4]~7 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[4]~7 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[5]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[5]~8 (
	.dataa(\av_ld_byte0_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_5),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[5]~8_combout ),
	.cout());
defparam \W_rf_wr_data[5]~8 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[5]~8 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[6]~9 (
	.dataa(\av_ld_byte0_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_6),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[6]~9_combout ),
	.cout());
defparam \W_rf_wr_data[6]~9 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[6]~9 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[7]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[1]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[7]~10 (
	.dataa(\av_ld_byte0_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_7),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[7]~10_combout ),
	.cout());
defparam \W_rf_wr_data[7]~10 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[7]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[8]~11 (
	.dataa(\av_ld_byte1_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_8),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[8]~11_combout ),
	.cout());
defparam \W_rf_wr_data[8]~11 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[8]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[9]~12 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_9),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[9]~12_combout ),
	.cout());
defparam \W_rf_wr_data[9]~12 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[9]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[10]~13 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_10),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[10]~13_combout ),
	.cout());
defparam \W_rf_wr_data[10]~13 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[10]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[11]~14 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_11),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[11]~14_combout ),
	.cout());
defparam \W_rf_wr_data[11]~14 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[11]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[12]~15 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_12),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[12]~15_combout ),
	.cout());
defparam \W_rf_wr_data[12]~15 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[12]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[13]~16 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_13),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[13]~16_combout ),
	.cout());
defparam \W_rf_wr_data[13]~16 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[13]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[14]~17 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_14),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[14]~17_combout ),
	.cout());
defparam \W_rf_wr_data[14]~17 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[14]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[15]~18 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_15),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[15]~18_combout ),
	.cout());
defparam \W_rf_wr_data[15]~18 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[15]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[16]~19 (
	.dataa(\av_ld_byte2_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_16),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[16]~19_combout ),
	.cout());
defparam \W_rf_wr_data[16]~19 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[16]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[17]~20 (
	.dataa(\av_ld_byte2_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_17),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[17]~20_combout ),
	.cout());
defparam \W_rf_wr_data[17]~20 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[17]~20 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[28]~21 (
	.dataa(\av_ld_byte3_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_28),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[28]~21_combout ),
	.cout());
defparam \W_rf_wr_data[28]~21 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[28]~21 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[27]~22 (
	.dataa(\av_ld_byte3_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_27),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[27]~22_combout ),
	.cout());
defparam \W_rf_wr_data[27]~22 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[27]~22 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[26]~23 (
	.dataa(\av_ld_byte3_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_26),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[26]~23_combout ),
	.cout());
defparam \W_rf_wr_data[26]~23 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[26]~23 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[25]~24 (
	.dataa(\av_ld_byte3_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_25),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[25]~24_combout ),
	.cout());
defparam \W_rf_wr_data[25]~24 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[25]~24 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[24]~25 (
	.dataa(\av_ld_byte3_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_24),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[24]~25_combout ),
	.cout());
defparam \W_rf_wr_data[24]~25 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[24]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[23]~26 (
	.dataa(\av_ld_byte2_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_23),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[23]~26_combout ),
	.cout());
defparam \W_rf_wr_data[23]~26 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[23]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[22]~27 (
	.dataa(\av_ld_byte2_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_22),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[22]~27_combout ),
	.cout());
defparam \W_rf_wr_data[22]~27 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[22]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[21]~28 (
	.dataa(\av_ld_byte2_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_21),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[21]~28_combout ),
	.cout());
defparam \W_rf_wr_data[21]~28 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[21]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[20]~29 (
	.dataa(\av_ld_byte2_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_20),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[20]~29_combout ),
	.cout());
defparam \W_rf_wr_data[20]~29 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[20]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[19]~30 (
	.dataa(\av_ld_byte2_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_19),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[19]~30_combout ),
	.cout());
defparam \W_rf_wr_data[19]~30 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[19]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[18]~31 (
	.dataa(\av_ld_byte2_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_18),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[18]~31_combout ),
	.cout());
defparam \W_rf_wr_data[18]~31 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[18]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~0 (
	.dataa(\Equal0~15_combout ),
	.datab(\Equal0~13_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.cout());
defparam \D_wr_dst_reg~0 .lut_mask = 16'hEFFF;
defparam \D_wr_dst_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~1 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\Equal0~16_combout ),
	.datac(\D_wr_dst_reg~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_wr_dst_reg~1_combout ),
	.cout());
defparam \D_wr_dst_reg~1 .lut_mask = 16'hFEFE;
defparam \D_wr_dst_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~17 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\Equal0~17_combout ),
	.cout());
defparam \Equal0~17 .lut_mask = 16'hAFFF;
defparam \Equal0~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 16'hFBFF;
defparam \D_ctrl_implicit_dst_eretaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~5 (
	.dataa(\D_iw[16]~q ),
	.datab(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~5_combout ),
	.cout());
defparam \D_dst_regnum[4]~5 .lut_mask = 16'hEEFF;
defparam \D_dst_regnum[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~6 (
	.dataa(\Equal62~9_combout ),
	.datab(\Equal62~14_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~6_combout ),
	.cout());
defparam \D_dst_regnum[4]~6 .lut_mask = 16'hEFFE;
defparam \D_dst_regnum[4]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~7 (
	.dataa(\Equal0~17_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\D_dst_regnum[4]~5_combout ),
	.datad(\D_dst_regnum[4]~6_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~7_combout ),
	.cout());
defparam \D_dst_regnum[4]~7 .lut_mask = 16'hFFFE;
defparam \D_dst_regnum[4]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~8 (
	.dataa(\D_dst_regnum[4]~7_combout ),
	.datab(\D_ctrl_exception~8_combout ),
	.datac(\D_ctrl_exception~14_combout ),
	.datad(\D_dst_regnum[4]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~8_combout ),
	.cout());
defparam \D_dst_regnum[4]~8 .lut_mask = 16'hBFFF;
defparam \D_dst_regnum[4]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~9 (
	.dataa(\D_dst_regnum[4]~8_combout ),
	.datab(\D_iw[26]~q ),
	.datac(\D_iw[21]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~9_combout ),
	.cout());
defparam \D_dst_regnum[4]~9 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[4]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~10 (
	.dataa(\D_dst_regnum[4]~8_combout ),
	.datab(\D_iw[22]~q ),
	.datac(\D_iw[17]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~10_combout ),
	.cout());
defparam \D_dst_regnum[0]~10 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[3]~11 (
	.dataa(\D_dst_regnum[4]~8_combout ),
	.datab(\D_iw[25]~q ),
	.datac(\D_iw[20]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~11_combout ),
	.cout());
defparam \D_dst_regnum[3]~11 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[3]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~12 (
	.dataa(\D_dst_regnum[4]~8_combout ),
	.datab(\D_iw[24]~q ),
	.datac(\D_iw[19]~q ),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~12_combout ),
	.cout());
defparam \D_dst_regnum[2]~12 .lut_mask = 16'hFAFC;
defparam \D_dst_regnum[2]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~18 (
	.dataa(\D_dst_regnum[4]~9_combout ),
	.datab(\D_dst_regnum[0]~10_combout ),
	.datac(\D_dst_regnum[3]~11_combout ),
	.datad(\D_dst_regnum[2]~12_combout ),
	.cin(gnd),
	.combout(\Equal0~18_combout ),
	.cout());
defparam \Equal0~18 .lut_mask = 16'h7FFF;
defparam \Equal0~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~13 (
	.dataa(\D_iw[23]~q ),
	.datab(\D_iw[18]~q ),
	.datac(gnd),
	.datad(\D_ctrl_b_is_dst~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~13_combout ),
	.cout());
defparam \D_dst_regnum[1]~13 .lut_mask = 16'hAACC;
defparam \D_dst_regnum[1]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~14 (
	.dataa(\Equal0~17_combout ),
	.datab(\D_dst_regnum[1]~13_combout ),
	.datac(gnd),
	.datad(\D_dst_regnum[4]~8_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~14_combout ),
	.cout());
defparam \D_dst_regnum[1]~14 .lut_mask = 16'hEEFF;
defparam \D_dst_regnum[1]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~2 (
	.dataa(\D_wr_dst_reg~1_combout ),
	.datab(\Equal0~18_combout ),
	.datac(gnd),
	.datad(\D_dst_regnum[1]~14_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~2_combout ),
	.cout());
defparam \D_wr_dst_reg~2 .lut_mask = 16'hFF77;
defparam \D_wr_dst_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~0 (
	.dataa(\W_alu_result[1]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.cout());
defparam \av_ld_rshift8~0 .lut_mask = 16'hEFFF;
defparam \av_ld_rshift8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~1 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_rshift8~1_combout ),
	.cout());
defparam \av_ld_rshift8~1 .lut_mask = 16'hEEEE;
defparam \av_ld_rshift8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data[1]~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\av_ld_rshift8~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data[1]~0_combout ),
	.cout());
defparam \av_ld_byte0_data[1]~0 .lut_mask = 16'hFF55;
defparam \av_ld_byte0_data[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(\D_iw[8]~q ),
	.datab(gnd),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.cout());
defparam \E_control_rd_data[0]~0 .lut_mask = 16'hAFFF;
defparam \E_control_rd_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~1 (
	.dataa(\D_iw[7]~q ),
	.datab(\W_estatus_reg~q ),
	.datac(\D_iw[6]~q ),
	.datad(\W_status_reg_pie~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~1_combout ),
	.cout());
defparam \E_control_rd_data[0]~1 .lut_mask = 16'hFFDE;
defparam \E_control_rd_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~2 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\D_iw[7]~q ),
	.datac(\E_control_rd_data[0]~1_combout ),
	.datad(\W_ienable_reg[0]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~2_combout ),
	.cout());
defparam \E_control_rd_data[0]~2 .lut_mask = 16'hFFBE;
defparam \E_control_rd_data[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~3 (
	.dataa(\W_ipending_reg[0]~q ),
	.datab(\E_control_rd_data[0]~0_combout ),
	.datac(\E_control_rd_data[0]~2_combout ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~3_combout ),
	.cout());
defparam \E_control_rd_data[0]~3 .lut_mask = 16'hFEFF;
defparam \E_control_rd_data[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~2 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(src_data_1),
	.datac(src_data_11),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~2_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~2 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[1]~4 (
	.dataa(\D_iw[7]~q ),
	.datab(\D_iw[6]~q ),
	.datac(\W_ienable_reg[1]~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[1]~4_combout ),
	.cout());
defparam \E_control_rd_data[1]~4 .lut_mask = 16'hFEFF;
defparam \E_control_rd_data[1]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[1]~5 (
	.dataa(\E_control_rd_data[1]~4_combout ),
	.datab(\W_ipending_reg[1]~q ),
	.datac(\E_control_rd_data[0]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_control_rd_data[1]~5_combout ),
	.cout());
defparam \E_control_rd_data[1]~5 .lut_mask = 16'hFEFE;
defparam \E_control_rd_data[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~3 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(src_data_2),
	.datac(src_data_21),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~3_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~3 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~4 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(src_data_3),
	.datac(src_data_31),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~4_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~4 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~5 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(src_data_4),
	.datac(src_data_41),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~5_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~5 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~6 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(src_data_5),
	.datac(src_data_51),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~6_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~6 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~7 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(src_data_6),
	.datac(src_data_61),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~7_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~7 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~8 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(src_data_7),
	.datac(src_data_71),
	.datad(\av_ld_rshift8~1_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~8_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~8 .lut_mask = 16'hFAFC;
defparam \av_ld_byte0_data_nxt[7]~8 .sum_lutc_input = "datac";

dffeas R_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_ld_signed~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cycloneive_lcell_comb \av_fill_bit~0 (
	.dataa(\R_ctrl_ld_signed~q ),
	.datab(\av_ld_byte1_data[7]~q ),
	.datac(\av_ld_byte0_data[7]~q ),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\av_fill_bit~0_combout ),
	.cout());
defparam \av_fill_bit~0 .lut_mask = 16'hFAFC;
defparam \av_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\D_ctrl_mem16~0_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.cout());
defparam \av_ld_byte1_data_en~0 .lut_mask = 16'hEFFF;
defparam \av_ld_byte1_data_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~0 (
	.dataa(out_data_buffer_282),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~0_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~0 .lut_mask = 16'hAFFA;
defparam \av_ld_byte3_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~1 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_28),
	.datad(out_data_buffer_283),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~1_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~1 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~2 (
	.dataa(src_payload6),
	.datab(\av_ld_byte3_data_nxt~1_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~2_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~2 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~3 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~0_combout ),
	.datac(\av_ld_byte3_data_nxt~2_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~3_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~3 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~4 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_27),
	.datad(av_readdata_pre_27),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~4_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~4 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~5 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_272),
	.datad(out_data_buffer_273),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~5_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~5 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~6 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~4_combout ),
	.datac(\av_ld_byte3_data_nxt~5_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~6_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~6 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~7 (
	.dataa(out_data_buffer_262),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~7_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~7 .lut_mask = 16'hAFFA;
defparam \av_ld_byte3_data_nxt~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~8 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_26),
	.datad(out_data_buffer_263),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~8_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~8 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~9 (
	.dataa(src_payload6),
	.datab(\av_ld_byte3_data_nxt~8_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~9_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~9 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~10 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~7_combout ),
	.datac(\av_ld_byte3_data_nxt~9_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~10_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~10 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~11 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_25),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~11_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~11 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~12 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_252),
	.datad(out_data_buffer_253),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~12_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~12 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~13 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~11_combout ),
	.datac(\av_ld_byte3_data_nxt~12_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~13_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~13 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~14 (
	.dataa(out_data_buffer_242),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~14_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~14 .lut_mask = 16'hAFFA;
defparam \av_ld_byte3_data_nxt~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~15 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_24),
	.datad(out_data_buffer_243),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~15_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~15 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~16 (
	.dataa(src_payload6),
	.datab(\av_ld_byte3_data_nxt~15_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~16_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~16 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~17 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~14_combout ),
	.datac(\av_ld_byte3_data_nxt~16_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~17_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~17 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~17 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

dffeas \av_ld_byte3_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

dffeas \av_ld_byte3_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[31]~32 (
	.dataa(\av_ld_byte3_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[31]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[31]~32_combout ),
	.cout());
defparam \W_rf_wr_data[31]~32 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[31]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[30]~33 (
	.dataa(\av_ld_byte3_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[30]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[30]~33_combout ),
	.cout());
defparam \W_rf_wr_data[30]~33 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[30]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[29]~34 (
	.dataa(\av_ld_byte3_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[29]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[29]~34_combout ),
	.cout());
defparam \W_rf_wr_data[29]~34 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[29]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~18 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_31),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~18_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~18 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~19 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_313),
	.datad(out_data_buffer_314),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~19_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~19 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~20 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~18_combout ),
	.datac(\av_ld_byte3_data_nxt~19_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~20_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~20 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~21 (
	.dataa(out_data_buffer_302),
	.datab(gnd),
	.datac(out_data_toggle_flopped),
	.datad(dreg_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~21_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~21 .lut_mask = 16'hAFFA;
defparam \av_ld_byte3_data_nxt~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~22 (
	.dataa(out_valid),
	.datab(src0_valid4),
	.datac(q_a_30),
	.datad(out_data_buffer_303),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~22_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~22 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~23 (
	.dataa(src_payload6),
	.datab(\av_ld_byte3_data_nxt~22_combout ),
	.datac(src0_valid2),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~23_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~23 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~24 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~21_combout ),
	.datac(\av_ld_byte3_data_nxt~23_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~24_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~24 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~25 (
	.dataa(src0_valid2),
	.datab(src0_valid4),
	.datac(q_a_29),
	.datad(av_readdata_pre_29),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~25_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~25 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~26 (
	.dataa(out_valid),
	.datab(out_valid1),
	.datac(out_data_buffer_292),
	.datad(out_data_buffer_293),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~26_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~26 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~27 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~25_combout ),
	.datac(\av_ld_byte3_data_nxt~26_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~27_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~27 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~9 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[0]~q ),
	.datad(src_data_0),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~9_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~9 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[0]~9 .sum_lutc_input = "datac";

dffeas \W_alu_result[28] (
	.clk(clk_clk),
	.d(\W_alu_result[28]~0_combout ),
	.asdata(\E_shift_rot_result[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_28),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \W_alu_result[27] (
	.clk(clk_clk),
	.d(\W_alu_result[27]~1_combout ),
	.asdata(\E_shift_rot_result[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_27),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(clk_clk),
	.d(\W_alu_result[26]~2_combout ),
	.asdata(\E_shift_rot_result[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_26),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(clk_clk),
	.d(\W_alu_result[25]~3_combout ),
	.asdata(\E_shift_rot_result[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_25),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(clk_clk),
	.d(\W_alu_result[24]~4_combout ),
	.asdata(\E_shift_rot_result[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_24),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(clk_clk),
	.d(\W_alu_result[23]~5_combout ),
	.asdata(\E_shift_rot_result[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_23),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(clk_clk),
	.d(\W_alu_result[22]~6_combout ),
	.asdata(\E_shift_rot_result[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_22),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(clk_clk),
	.d(\W_alu_result[21]~7_combout ),
	.asdata(\E_shift_rot_result[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_21),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(clk_clk),
	.d(\W_alu_result[20]~8_combout ),
	.asdata(\E_shift_rot_result[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_20),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(clk_clk),
	.d(\W_alu_result[19]~9_combout ),
	.asdata(\E_shift_rot_result[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_19),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(clk_clk),
	.d(\W_alu_result[18]~10_combout ),
	.asdata(\E_shift_rot_result[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_18),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(clk_clk),
	.d(\W_alu_result[17]~11_combout ),
	.asdata(\E_shift_rot_result[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_17),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(clk_clk),
	.d(\W_alu_result[16]~12_combout ),
	.asdata(\E_shift_rot_result[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_16),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(clk_clk),
	.d(\W_alu_result[15]~13_combout ),
	.asdata(\E_shift_rot_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(clk_clk),
	.d(\W_alu_result[14]~14_combout ),
	.asdata(\E_shift_rot_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(clk_clk),
	.d(\W_alu_result[13]~15_combout ),
	.asdata(\E_shift_rot_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[6] (
	.clk(clk_clk),
	.d(\W_alu_result[6]~22_combout ),
	.asdata(\E_shift_rot_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[7] (
	.clk(clk_clk),
	.d(\W_alu_result[7]~21_combout ),
	.asdata(\E_shift_rot_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(clk_clk),
	.d(\W_alu_result[5]~23_combout ),
	.asdata(\E_shift_rot_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[4] (
	.clk(clk_clk),
	.d(\W_alu_result[4]~24_combout ),
	.asdata(\E_shift_rot_result[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[12] (
	.clk(clk_clk),
	.d(\W_alu_result[12]~16_combout ),
	.asdata(\E_shift_rot_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(clk_clk),
	.d(\W_alu_result[10]~18_combout ),
	.asdata(\E_shift_rot_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(clk_clk),
	.d(\W_alu_result[9]~19_combout ),
	.asdata(\E_shift_rot_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(clk_clk),
	.d(\W_alu_result[8]~20_combout ),
	.asdata(\E_shift_rot_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(clk_clk),
	.d(\W_alu_result[11]~17_combout ),
	.asdata(\E_shift_rot_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(clk_clk),
	.d(\W_alu_result[2]~25_combout ),
	.asdata(\E_shift_rot_result[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(clk_clk),
	.d(\W_alu_result[3]~26_combout ),
	.asdata(\E_shift_rot_result[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\d_writedata[31]~3_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\d_writedata[30]~4_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\d_writedata[29]~5_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\d_writedata[28]~6_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\d_writedata[27]~7_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\d_writedata[26]~2_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\d_writedata[25]~1_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\d_writedata[24]~0_combout ),
	.asdata(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \F_pc[26] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[26]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_26),
	.prn(vcc));
defparam \F_pc[26] .is_wysiwyg = "true";
defparam \F_pc[26] .power_up = "low";

dffeas \F_pc[25] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[25]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_25),
	.prn(vcc));
defparam \F_pc[25] .is_wysiwyg = "true";
defparam \F_pc[25] .power_up = "low";

dffeas \F_pc[24] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[24]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_24),
	.prn(vcc));
defparam \F_pc[24] .is_wysiwyg = "true";
defparam \F_pc[24] .power_up = "low";

dffeas \F_pc[23] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[23]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_23),
	.prn(vcc));
defparam \F_pc[23] .is_wysiwyg = "true";
defparam \F_pc[23] .power_up = "low";

dffeas \F_pc[22] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[22]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_22),
	.prn(vcc));
defparam \F_pc[22] .is_wysiwyg = "true";
defparam \F_pc[22] .power_up = "low";

dffeas \F_pc[21] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[21]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_21),
	.prn(vcc));
defparam \F_pc[21] .is_wysiwyg = "true";
defparam \F_pc[21] .power_up = "low";

dffeas \F_pc[20] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[20]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_20),
	.prn(vcc));
defparam \F_pc[20] .is_wysiwyg = "true";
defparam \F_pc[20] .power_up = "low";

dffeas \F_pc[19] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[19]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_19),
	.prn(vcc));
defparam \F_pc[19] .is_wysiwyg = "true";
defparam \F_pc[19] .power_up = "low";

dffeas \F_pc[18] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[18]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_18),
	.prn(vcc));
defparam \F_pc[18] .is_wysiwyg = "true";
defparam \F_pc[18] .power_up = "low";

dffeas \F_pc[17] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[17]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_17),
	.prn(vcc));
defparam \F_pc[17] .is_wysiwyg = "true";
defparam \F_pc[17] .power_up = "low";

dffeas \F_pc[16] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[16]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_16),
	.prn(vcc));
defparam \F_pc[16] .is_wysiwyg = "true";
defparam \F_pc[16] .power_up = "low";

dffeas \F_pc[15] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[15]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_15),
	.prn(vcc));
defparam \F_pc[15] .is_wysiwyg = "true";
defparam \F_pc[15] .power_up = "low";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[14]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_14),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[13]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[12]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[11]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[10]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[8]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[7]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[6]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[5]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[3]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[2]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[4]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[9]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[0]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[1]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\E_st_data[8]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\E_st_data[9]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\E_st_data[10]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\E_st_data[11]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\E_st_data[12]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\E_st_data[13]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\E_st_data[14]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\E_st_data[15]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\E_st_data[16]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\E_st_data[17]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\E_st_data[21]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\E_st_data[18]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\E_st_data[23]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\E_st_data[22]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\E_st_data[20]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\E_st_data[19]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

cycloneive_lcell_comb \av_ld_getting_data~9 (
	.dataa(read_latency_shift_reg_02),
	.datab(mem_67_07),
	.datac(WideOr1),
	.datad(\av_ld_getting_data~7_combout ),
	.cin(gnd),
	.combout(av_ld_getting_data),
	.cout());
defparam \av_ld_getting_data~9 .lut_mask = 16'hFFF7;
defparam \av_ld_getting_data~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_valid~0 (
	.dataa(av_readdatavalid),
	.datab(gnd),
	.datac(gnd),
	.datad(i_read1),
	.cin(gnd),
	.combout(\F_valid~0_combout ),
	.cout());
defparam \F_valid~0 .lut_mask = 16'hAAFF;
defparam \F_valid~0 .sum_lutc_input = "datac";

dffeas D_valid(
	.clk(clk_clk),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(clk_clk),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

cycloneive_lcell_comb \av_ld_getting_data~2 (
	.dataa(mem_67_0),
	.datab(src0_valid),
	.datac(mem_67_01),
	.datad(src0_valid1),
	.cin(gnd),
	.combout(\av_ld_getting_data~2_combout ),
	.cout());
defparam \av_ld_getting_data~2 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~3 (
	.dataa(mem_67_02),
	.datab(src0_valid2),
	.datac(mem_67_03),
	.datad(src0_valid3),
	.cin(gnd),
	.combout(\av_ld_getting_data~3_combout ),
	.cout());
defparam \av_ld_getting_data~3 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~4 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_67_04),
	.datac(read_latency_shift_reg_03),
	.datad(mem_67_05),
	.cin(gnd),
	.combout(\av_ld_getting_data~4_combout ),
	.cout());
defparam \av_ld_getting_data~4 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~5 (
	.dataa(\av_ld_getting_data~4_combout ),
	.datab(gnd),
	.datac(mem_67_06),
	.datad(src0_valid4),
	.cin(gnd),
	.combout(\av_ld_getting_data~5_combout ),
	.cout());
defparam \av_ld_getting_data~5 .lut_mask = 16'hAFFF;
defparam \av_ld_getting_data~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~6 (
	.dataa(out_valid),
	.datab(out_data_buffer_67),
	.datac(out_valid1),
	.datad(out_data_buffer_671),
	.cin(gnd),
	.combout(\av_ld_getting_data~6_combout ),
	.cout());
defparam \av_ld_getting_data~6 .lut_mask = 16'h7FFF;
defparam \av_ld_getting_data~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~7 (
	.dataa(\av_ld_getting_data~2_combout ),
	.datab(\av_ld_getting_data~3_combout ),
	.datac(\av_ld_getting_data~5_combout ),
	.datad(\av_ld_getting_data~6_combout ),
	.cin(gnd),
	.combout(\av_ld_getting_data~7_combout ),
	.cout());
defparam \av_ld_getting_data~7 .lut_mask = 16'hFFFE;
defparam \av_ld_getting_data~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_getting_data~8 (
	.dataa(src_payload),
	.datab(d_read1),
	.datac(WideOr1),
	.datad(\av_ld_getting_data~7_combout ),
	.cin(gnd),
	.combout(\av_ld_getting_data~8_combout ),
	.cout());
defparam \av_ld_getting_data~8 .lut_mask = 16'hBFFF;
defparam \av_ld_getting_data~8 .sum_lutc_input = "datac";

dffeas E_new_inst(
	.clk(clk_clk),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

cycloneive_lcell_comb \F_iw[2]~13 (
	.dataa(src_payload3),
	.datab(src1_valid),
	.datac(readdata_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[2]~13_combout ),
	.cout());
defparam \F_iw[2]~13 .lut_mask = 16'hFEFE;
defparam \F_iw[2]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~14 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_2),
	.datad(av_readdata_pre_2),
	.cin(gnd),
	.combout(\F_iw[2]~14_combout ),
	.cout());
defparam \F_iw[2]~14 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~15 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_2),
	.datad(out_data_buffer_21),
	.cin(gnd),
	.combout(\F_iw[2]~15_combout ),
	.cout());
defparam \F_iw[2]~15 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~16 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[2]~13_combout ),
	.datac(\F_iw[2]~14_combout ),
	.datad(\F_iw[2]~15_combout ),
	.cin(gnd),
	.combout(\F_iw[2]~16_combout ),
	.cout());
defparam \F_iw[2]~16 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~16 .sum_lutc_input = "datac";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

cycloneive_lcell_comb \F_iw[0]~4 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_0),
	.datad(av_readdata_pre_0),
	.cin(gnd),
	.combout(\F_iw[0]~4_combout ),
	.cout());
defparam \F_iw[0]~4 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~5 (
	.dataa(src_payload3),
	.datab(\F_iw[0]~4_combout ),
	.datac(src1_valid),
	.datad(readdata_0),
	.cin(gnd),
	.combout(\F_iw[0]~5_combout ),
	.cout());
defparam \F_iw[0]~5 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~6 (
	.dataa(read_latency_shift_reg_04),
	.datab(mem_86_01),
	.datac(mem_68_01),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(\F_iw[0]~6_combout ),
	.cout());
defparam \F_iw[0]~6 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~7 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_0),
	.datad(out_data_buffer_01),
	.cin(gnd),
	.combout(\F_iw[0]~7_combout ),
	.cout());
defparam \F_iw[0]~7 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~8 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[0]~5_combout ),
	.datac(\F_iw[0]~6_combout ),
	.datad(\F_iw[0]~7_combout ),
	.cin(gnd),
	.combout(\F_iw[0]~8_combout ),
	.cout());
defparam \F_iw[0]~8 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~8 .sum_lutc_input = "datac";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cycloneive_lcell_comb \F_iw[1]~9 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_1),
	.datad(av_readdata_pre_1),
	.cin(gnd),
	.combout(\F_iw[1]~9_combout ),
	.cout());
defparam \F_iw[1]~9 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[1]~10 (
	.dataa(src_payload1),
	.datab(out_valid2),
	.datac(out_data_buffer_1),
	.datad(av_readdata_pre_11),
	.cin(gnd),
	.combout(\F_iw[1]~10_combout ),
	.cout());
defparam \F_iw[1]~10 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[1]~11 (
	.dataa(\F_iw[1]~9_combout ),
	.datab(\F_iw[1]~10_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_11),
	.cin(gnd),
	.combout(\F_iw[1]~11_combout ),
	.cout());
defparam \F_iw[1]~11 .lut_mask = 16'hFFFE;
defparam \F_iw[1]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[1]~12 (
	.dataa(\F_iw[1]~11_combout ),
	.datab(src1_valid),
	.datac(readdata_1),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[1]~12_combout ),
	.cout());
defparam \F_iw[1]~12 .lut_mask = 16'hFEFF;
defparam \F_iw[1]~12 .sum_lutc_input = "datac";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cycloneive_lcell_comb \F_iw[4]~21 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_4),
	.datad(readdata_4),
	.cin(gnd),
	.combout(\F_iw[4]~21_combout ),
	.cout());
defparam \F_iw[4]~21 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[4]~22 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_4),
	.datad(q_a_4),
	.cin(gnd),
	.combout(\F_iw[4]~22_combout ),
	.cout());
defparam \F_iw[4]~22 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[4]~23 (
	.dataa(\F_iw[4]~21_combout ),
	.datab(\F_iw[4]~22_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_41),
	.cin(gnd),
	.combout(\F_iw[4]~23_combout ),
	.cout());
defparam \F_iw[4]~23 .lut_mask = 16'hFFFE;
defparam \F_iw[4]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[4]~24 (
	.dataa(src_payload3),
	.datab(\F_iw[4]~23_combout ),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[4]~24_combout ),
	.cout());
defparam \F_iw[4]~24 .lut_mask = 16'hEEFF;
defparam \F_iw[4]~24 .sum_lutc_input = "datac";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cycloneive_lcell_comb \F_iw[3]~17 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_3),
	.datad(readdata_31),
	.cin(gnd),
	.combout(\F_iw[3]~17_combout ),
	.cout());
defparam \F_iw[3]~17 .lut_mask = 16'hFFFE;
defparam \F_iw[3]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[3]~18 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_3),
	.datad(q_a_3),
	.cin(gnd),
	.combout(\F_iw[3]~18_combout ),
	.cout());
defparam \F_iw[3]~18 .lut_mask = 16'hFFFE;
defparam \F_iw[3]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[3]~19 (
	.dataa(\F_iw[3]~17_combout ),
	.datab(\F_iw[3]~18_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_31),
	.cin(gnd),
	.combout(\F_iw[3]~19_combout ),
	.cout());
defparam \F_iw[3]~19 .lut_mask = 16'hFFFE;
defparam \F_iw[3]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[3]~20 (
	.dataa(src_payload3),
	.datab(\F_iw[3]~19_combout ),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[3]~20_combout ),
	.cout());
defparam \F_iw[3]~20 .lut_mask = 16'hEEFF;
defparam \F_iw[3]~20 .sum_lutc_input = "datac";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.cout());
defparam \D_ctrl_ld_signed~0 .lut_mask = 16'hEFFF;
defparam \D_ctrl_ld_signed~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld~2_combout ),
	.cout());
defparam \D_ctrl_ld~2 .lut_mask = 16'hBFBF;
defparam \D_ctrl_ld~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~3 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(\D_iw[0]~q ),
	.datad(\D_ctrl_ld~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_ld~3_combout ),
	.cout());
defparam \D_ctrl_ld~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_ld~3 .sum_lutc_input = "datac";

dffeas R_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

dffeas av_ld_waiting_for_data(
	.clk(clk_clk),
	.d(\av_ld_waiting_for_data_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cycloneive_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(\av_ld_getting_data~8_combout ),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_ld~q ),
	.datad(\av_ld_waiting_for_data~q ),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 16'hFAFC;
defparam \av_ld_waiting_for_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFBFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~37 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_5),
	.datad(av_readdata_pre_5),
	.cin(gnd),
	.combout(\F_iw[5]~37_combout ),
	.cout());
defparam \F_iw[5]~37 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~38 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_5),
	.datad(out_data_buffer_51),
	.cin(gnd),
	.combout(\F_iw[5]~38_combout ),
	.cout());
defparam \F_iw[5]~38 .lut_mask = 16'hFFFE;
defparam \F_iw[5]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~39 (
	.dataa(src_payload5),
	.datab(\F_iw[5]~37_combout ),
	.datac(\F_iw[5]~38_combout ),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[5]~39_combout ),
	.cout());
defparam \F_iw[5]~39 .lut_mask = 16'hFEFF;
defparam \F_iw[5]~39 .sum_lutc_input = "datac";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cycloneive_lcell_comb \Equal0~7 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~2_combout ),
	.datac(\D_iw[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'hFEFE;
defparam \Equal0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~43 (
	.dataa(src1_valid1),
	.datab(av_readdata_pre_15),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[15]~43_combout ),
	.cout());
defparam \F_iw[15]~43 .lut_mask = 16'hEEFF;
defparam \F_iw[15]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~44 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_15),
	.datad(out_data_buffer_151),
	.cin(gnd),
	.combout(\F_iw[15]~44_combout ),
	.cout());
defparam \F_iw[15]~44 .lut_mask = 16'hFFFE;
defparam \F_iw[15]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~45 (
	.dataa(\F_iw[15]~43_combout ),
	.datab(\F_iw[15]~44_combout ),
	.datac(src1_valid2),
	.datad(q_a_15),
	.cin(gnd),
	.combout(\F_iw[15]~45_combout ),
	.cout());
defparam \F_iw[15]~45 .lut_mask = 16'hFFFE;
defparam \F_iw[15]~45 .sum_lutc_input = "datac";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_st~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.cout());
defparam \D_ctrl_st~0 .lut_mask = 16'hBFFF;
defparam \D_ctrl_st~0 .sum_lutc_input = "datac";

dffeas R_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cycloneive_lcell_comb \W_valid~3 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\E_valid_from_R~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_valid~3_combout ),
	.cout());
defparam \W_valid~3 .lut_mask = 16'hF7F7;
defparam \W_valid~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_valid~2 (
	.dataa(\E_stall~4_combout ),
	.datab(d_write1),
	.datac(av_waitrequest),
	.datad(\W_valid~3_combout ),
	.cin(gnd),
	.combout(\W_valid~2_combout ),
	.cout());
defparam \W_valid~2 .lut_mask = 16'hFF7F;
defparam \W_valid~2 .sum_lutc_input = "datac";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cycloneive_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(\hbreak_pending~q ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.cout());
defparam \hbreak_pending_nxt~0 .lut_mask = 16'hEEFF;
defparam \hbreak_pending_nxt~0 .sum_lutc_input = "datac";

dffeas hbreak_pending(
	.clk(clk_clk),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cycloneive_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datab(hbreak_enabled1),
	.datac(\wait_for_one_post_bret_inst~q ),
	.datad(\F_valid~0_combout ),
	.cin(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.cout());
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 16'hFEFF;
defparam \wait_for_one_post_bret_inst~0 .sum_lutc_input = "datac";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cycloneive_lcell_comb \hbreak_req~0 (
	.dataa(\W_valid~q ),
	.datab(\hbreak_pending~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|jtag_break~q ),
	.datad(\wait_for_one_post_bret_inst~q ),
	.cin(gnd),
	.combout(\hbreak_req~0_combout ),
	.cout());
defparam \hbreak_req~0 .lut_mask = 16'hFEFF;
defparam \hbreak_req~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~40 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_14),
	.datad(q_a_14),
	.cin(gnd),
	.combout(\F_iw[14]~40_combout ),
	.cout());
defparam \F_iw[14]~40 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~41 (
	.dataa(src_payload3),
	.datab(\F_iw[14]~40_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\F_iw[14]~41_combout ),
	.cout());
defparam \F_iw[14]~41 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~42 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[14]~41_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_141),
	.cin(gnd),
	.combout(\F_iw[14]~42_combout ),
	.cout());
defparam \F_iw[14]~42 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~110 (
	.dataa(\D_iw[26]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[14]~42_combout ),
	.cin(gnd),
	.combout(\F_iw[14]~110_combout ),
	.cout());
defparam \F_iw[14]~110 .lut_mask = 16'hFFDF;
defparam \F_iw[14]~110 .sum_lutc_input = "datac";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~110_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cycloneive_lcell_comb \D_op_opx_rsv63~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_op_opx_rsv63~0_combout ),
	.cout());
defparam \D_op_opx_rsv63~0 .lut_mask = 16'hEEEE;
defparam \D_op_opx_rsv63~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~28 (
	.dataa(src1_valid1),
	.datab(av_readdata_pre_13),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[13]~28_combout ),
	.cout());
defparam \F_iw[13]~28 .lut_mask = 16'hEEFF;
defparam \F_iw[13]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~29 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_13),
	.datad(out_data_buffer_131),
	.cin(gnd),
	.combout(\F_iw[13]~29_combout ),
	.cout());
defparam \F_iw[13]~29 .lut_mask = 16'hFFFE;
defparam \F_iw[13]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~30 (
	.dataa(\F_iw[13]~28_combout ),
	.datab(\F_iw[13]~29_combout ),
	.datac(src1_valid2),
	.datad(q_a_13),
	.cin(gnd),
	.combout(\F_iw[13]~30_combout ),
	.cout());
defparam \F_iw[13]~30 .lut_mask = 16'hFFFE;
defparam \F_iw[13]~30 .sum_lutc_input = "datac";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

cycloneive_lcell_comb \F_iw[16]~31 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_16),
	.datad(av_readdata_pre_16),
	.cin(gnd),
	.combout(\F_iw[16]~31_combout ),
	.cout());
defparam \F_iw[16]~31 .lut_mask = 16'hFFFE;
defparam \F_iw[16]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[16]~32 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_16),
	.datad(out_data_buffer_161),
	.cin(gnd),
	.combout(\F_iw[16]~32_combout ),
	.cout());
defparam \F_iw[16]~32 .lut_mask = 16'hFFFE;
defparam \F_iw[16]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[16]~33 (
	.dataa(src_payload4),
	.datab(\F_iw[16]~31_combout ),
	.datac(\F_iw[16]~32_combout ),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[16]~33_combout ),
	.cout());
defparam \F_iw[16]~33 .lut_mask = 16'hFEFF;
defparam \F_iw[16]~33 .sum_lutc_input = "datac";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cycloneive_lcell_comb \F_iw[12]~34 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_12),
	.datad(av_readdata_pre_12),
	.cin(gnd),
	.combout(\F_iw[12]~34_combout ),
	.cout());
defparam \F_iw[12]~34 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[12]~35 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_12),
	.datad(out_data_buffer_121),
	.cin(gnd),
	.combout(\F_iw[12]~35_combout ),
	.cout());
defparam \F_iw[12]~35 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[12]~36 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[12]~34_combout ),
	.datac(\F_iw[12]~35_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[12]~36_combout ),
	.cout());
defparam \F_iw[12]~36 .lut_mask = 16'hFEFE;
defparam \F_iw[12]~36 .sum_lutc_input = "datac";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~36_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cycloneive_lcell_comb \Equal62~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~4_combout ),
	.cout());
defparam \Equal62~4 .lut_mask = 16'hFF7F;
defparam \Equal62~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~5 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~5_combout ),
	.cout());
defparam \Equal62~5 .lut_mask = 16'hFFF7;
defparam \Equal62~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~6 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~6_combout ),
	.cout());
defparam \Equal62~6 .lut_mask = 16'hFFFB;
defparam \Equal62~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~5_combout ),
	.datad(\Equal62~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~7 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~7_combout ),
	.cout());
defparam \Equal62~7 .lut_mask = 16'hFFBF;
defparam \Equal62~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(\Equal62~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_shift_rot~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(\D_iw[12]~q ),
	.datab(gnd),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.cout());
defparam \D_ctrl_shift_logical~0 .lut_mask = 16'hAFFF;
defparam \D_ctrl_shift_logical~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.cout());
defparam \D_ctrl_shift_rot~2 .lut_mask = 16'hACFF;
defparam \D_ctrl_shift_rot~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~3 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_shift_rot~0_combout ),
	.datac(\D_ctrl_shift_rot~1_combout ),
	.datad(\D_ctrl_shift_rot~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~3_combout ),
	.cout());
defparam \D_ctrl_shift_rot~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~3 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[0]~5 (
	.dataa(\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\E_shift_rot_cnt[0]~5_combout ),
	.cout(\E_shift_rot_cnt[0]~6 ));
defparam \E_shift_rot_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \E_shift_rot_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~0 .lut_mask = 16'hFFF7;
defparam \D_ctrl_hi_imm16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\D_ctrl_hi_imm16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~1_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~1 .lut_mask = 16'hFEFE;
defparam \D_ctrl_hi_imm16~1 .sum_lutc_input = "datac";

dffeas R_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_hi_imm16~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[0]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~14_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~14 .lut_mask = 16'hF6FF;
defparam \D_ctrl_alu_force_xor~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~14_combout ),
	.cout());
defparam \Equal0~14 .lut_mask = 16'hFFFE;
defparam \Equal0~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~15 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~15_combout ),
	.cout());
defparam \Equal0~15 .lut_mask = 16'hFFFD;
defparam \Equal0~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_ctrl_alu_force_xor~14_combout ),
	.datac(\Equal0~14_combout ),
	.datad(\Equal0~15_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~3_combout ),
	.cout());
defparam \D_dst_regnum[4]~3 .lut_mask = 16'h7FFF;
defparam \D_dst_regnum[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~8 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~8_combout ),
	.cout());
defparam \Equal62~8 .lut_mask = 16'hFEFF;
defparam \Equal62~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~14 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~14_combout ),
	.cout());
defparam \Equal62~14 .lut_mask = 16'hFDFF;
defparam \Equal62~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~8_combout ),
	.datac(\Equal62~14_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~12 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~12_combout ),
	.cout());
defparam \Equal62~12 .lut_mask = 16'hEFFF;
defparam \Equal62~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal62~12_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~10_combout ),
	.cout());
defparam \Equal62~10 .lut_mask = 16'hBFFF;
defparam \Equal62~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(\D_iw[15]~q ),
	.datab(gnd),
	.datac(\Equal0~7_combout ),
	.datad(\Equal62~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 16'hAFFF;
defparam \D_ctrl_uncond_cti_non_br~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~13 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~13_combout ),
	.cout());
defparam \Equal0~13 .lut_mask = 16'hDFFF;
defparam \Equal0~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~9 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~9_combout ),
	.cout());
defparam \Equal62~9 .lut_mask = 16'hFFEF;
defparam \Equal62~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hEEEE;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_cmpge~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_cmpge~0_combout ),
	.cout());
defparam \D_op_cmpge~0 .lut_mask = 16'hFEFF;
defparam \D_op_cmpge~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~4 (
	.dataa(gnd),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~4_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~4_combout ),
	.cout());
defparam \D_ctrl_exception~4 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~11 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~11_combout ),
	.cout());
defparam \Equal62~11 .lut_mask = 16'hDFFF;
defparam \Equal62~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv17~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv17~0_combout ),
	.cout());
defparam \D_op_opx_rsv17~0 .lut_mask = 16'hFEFF;
defparam \D_op_opx_rsv17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~5 (
	.dataa(gnd),
	.datab(\Equal62~10_combout ),
	.datac(\Equal62~11_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~5_combout ),
	.cout());
defparam \D_ctrl_exception~5 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~2_combout ),
	.cout());
defparam \Equal62~2 .lut_mask = 16'hFBFF;
defparam \Equal62~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv00~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv00~0_combout ),
	.cout());
defparam \D_op_opx_rsv00~0 .lut_mask = 16'hEFFF;
defparam \D_op_opx_rsv00~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~6 (
	.dataa(gnd),
	.datab(\Equal62~2_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~6_combout ),
	.cout());
defparam \D_ctrl_exception~6 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~7 (
	.dataa(gnd),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~6_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~7_combout ),
	.cout());
defparam \D_ctrl_exception~7 .lut_mask = 16'h3FFF;
defparam \D_ctrl_exception~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~8 (
	.dataa(\D_ctrl_exception~4_combout ),
	.datab(\D_ctrl_exception~5_combout ),
	.datac(\D_ctrl_exception~6_combout ),
	.datad(\D_ctrl_exception~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~8_combout ),
	.cout());
defparam \D_ctrl_exception~8 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~11 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~11_combout ),
	.cout());
defparam \Equal0~11 .lut_mask = 16'hFDFF;
defparam \Equal0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~9 (
	.dataa(\Equal62~6_combout ),
	.datab(\Equal62~5_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_exception~9_combout ),
	.cout());
defparam \D_ctrl_exception~9 .lut_mask = 16'h7F7F;
defparam \D_ctrl_exception~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~10 (
	.dataa(\D_op_opx_rsv17~0_combout ),
	.datab(\Equal62~6_combout ),
	.datac(\Equal62~5_combout ),
	.datad(\Equal62~12_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~10_combout ),
	.cout());
defparam \D_ctrl_exception~10 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~13 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~13_combout ),
	.cout());
defparam \Equal62~13 .lut_mask = 16'hFFFE;
defparam \Equal62~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~11 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_exception~11_combout ),
	.cout());
defparam \D_ctrl_exception~11 .lut_mask = 16'h7F7F;
defparam \D_ctrl_exception~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~3 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~3_combout ),
	.cout());
defparam \Equal62~3 .lut_mask = 16'hFFFD;
defparam \Equal62~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~1_combout ),
	.cout());
defparam \Equal62~1 .lut_mask = 16'hF7FF;
defparam \Equal62~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~12 (
	.dataa(\Equal62~14_combout ),
	.datab(\Equal62~3_combout ),
	.datac(\Equal62~1_combout ),
	.datad(\Equal62~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~12_combout ),
	.cout());
defparam \D_ctrl_exception~12 .lut_mask = 16'h7FFF;
defparam \D_ctrl_exception~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~13 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_op_opx_rsv63~0_combout ),
	.datac(\D_ctrl_exception~11_combout ),
	.datad(\D_ctrl_exception~12_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~13_combout ),
	.cout());
defparam \D_ctrl_exception~13 .lut_mask = 16'hFFF7;
defparam \D_ctrl_exception~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~14 (
	.dataa(\Equal0~11_combout ),
	.datab(\D_ctrl_exception~9_combout ),
	.datac(\D_ctrl_exception~10_combout ),
	.datad(\D_ctrl_exception~13_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~14_combout ),
	.cout());
defparam \D_ctrl_exception~14 .lut_mask = 16'hFFFD;
defparam \D_ctrl_exception~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~11_combout ),
	.datac(\Equal62~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.cout());
defparam \D_ctrl_retaddr~0 .lut_mask = 16'hFEFE;
defparam \D_ctrl_retaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(\Equal62~8_combout ),
	.datab(\Equal62~14_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.cout());
defparam \D_ctrl_retaddr~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_retaddr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_retaddr~0_combout ),
	.datad(\D_ctrl_retaddr~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.cout());
defparam \D_ctrl_retaddr~2 .lut_mask = 16'hFFFE;
defparam \D_ctrl_retaddr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'h7FFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~12 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~12_combout ),
	.cout());
defparam \Equal0~12 .lut_mask = 16'hBFFF;
defparam \Equal0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~12_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.cout());
defparam \D_ctrl_retaddr~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_retaddr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~2_combout ),
	.datac(\D_ctrl_retaddr~2_combout ),
	.datad(\D_ctrl_retaddr~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 16'hBFFF;
defparam \D_ctrl_force_src2_zero~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~3 (
	.dataa(\D_ctrl_exception~8_combout ),
	.datab(\D_ctrl_exception~14_combout ),
	.datac(\D_ctrl_force_src2_zero~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~3_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_force_src2_zero~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~4 (
	.dataa(\D_ctrl_force_src2_zero~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~1_combout ),
	.datac(\Equal0~13_combout ),
	.datad(\D_ctrl_force_src2_zero~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~4_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~4 .lut_mask = 16'hFFDF;
defparam \D_ctrl_force_src2_zero~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~5 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~12_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~5_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~5 .lut_mask = 16'hFFDE;
defparam \D_ctrl_force_src2_zero~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~6 (
	.dataa(\D_dst_regnum[4]~3_combout ),
	.datab(\D_ctrl_force_src2_zero~4_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_force_src2_zero~5_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~6_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~6 .lut_mask = 16'hFFF7;
defparam \D_ctrl_force_src2_zero~6 .sum_lutc_input = "datac";

dffeas R_ctrl_force_src2_zero(
	.clk(clk_clk),
	.d(\D_ctrl_force_src2_zero~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

cycloneive_lcell_comb \R_src2_lo[4]~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\R_ctrl_hi_imm16~q ),
	.datad(\R_ctrl_force_src2_zero~q ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~11_combout ),
	.cout());
defparam \R_src2_lo[4]~11 .lut_mask = 16'h0FFF;
defparam \R_src2_lo[4]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~100 (
	.dataa(src1_valid),
	.datab(src_payload2),
	.datac(av_readdata_pre_30),
	.datad(readdata_6),
	.cin(gnd),
	.combout(\F_iw[6]~100_combout ),
	.cout());
defparam \F_iw[6]~100 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~101 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_6),
	.datad(av_readdata_pre_6),
	.cin(gnd),
	.combout(\F_iw[6]~101_combout ),
	.cout());
defparam \F_iw[6]~101 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~101 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~102 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_6),
	.datad(out_data_buffer_61),
	.cin(gnd),
	.combout(\F_iw[6]~102_combout ),
	.cout());
defparam \F_iw[6]~102 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~102 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~103 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[6]~100_combout ),
	.datac(\F_iw[6]~101_combout ),
	.datad(\F_iw[6]~102_combout ),
	.cin(gnd),
	.combout(\F_iw[6]~103_combout ),
	.cout());
defparam \F_iw[6]~103 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~103 .sum_lutc_input = "datac";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~103_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cycloneive_lcell_comb \D_dst_regnum[4]~0 (
	.dataa(\D_iw[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~0_combout ),
	.cout());
defparam \D_dst_regnum[4]~0 .lut_mask = 16'hAAFF;
defparam \D_dst_regnum[4]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~2 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~4_combout ),
	.datad(\D_dst_regnum[4]~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_unsigned_lo_imm16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~5 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~2_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_unsigned_lo_imm16~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~16 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~16_combout ),
	.cout());
defparam \Equal0~16 .lut_mask = 16'hFFDF;
defparam \Equal0~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~0 .lut_mask = 16'h6996;
defparam \D_ctrl_b_is_dst~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~1_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~1 .lut_mask = 16'hFBFE;
defparam \D_ctrl_b_is_dst~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~2 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_ctrl_b_is_dst~0_combout ),
	.datad(\D_ctrl_b_is_dst~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~2_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~2 .lut_mask = 16'h96FF;
defparam \D_ctrl_b_is_dst~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~0 (
	.dataa(\Equal0~16_combout ),
	.datab(\D_ctrl_b_is_dst~2_combout ),
	.datac(\Equal0~15_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.cout());
defparam \R_src2_use_imm~0 .lut_mask = 16'hFEFF;
defparam \R_src2_use_imm~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.cout());
defparam \R_ctrl_br_nxt~0 .lut_mask = 16'hFFFE;
defparam \R_ctrl_br_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~1 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~1_combout ),
	.cout());
defparam \R_ctrl_br_nxt~1 .lut_mask = 16'hEEFF;
defparam \R_ctrl_br_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~1 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\R_src2_use_imm~0_combout ),
	.datac(\R_valid~q ),
	.datad(\R_ctrl_br_nxt~1_combout ),
	.cin(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.cout());
defparam \R_src2_use_imm~1 .lut_mask = 16'hFFFE;
defparam \R_src2_use_imm~1 .sum_lutc_input = "datac";

dffeas R_src2_use_imm(
	.clk(clk_clk),
	.d(\R_src2_use_imm~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 16'hBBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 16'hEFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .sum_lutc_input = "datac";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cycloneive_lcell_comb \E_src2[0]~16 (
	.dataa(\R_src2_use_imm~q ),
	.datab(\R_ctrl_src_imm5_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[0]~16_combout ),
	.cout());
defparam \E_src2[0]~16 .lut_mask = 16'hEEEE;
defparam \E_src2[0]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[0]~16 (
	.dataa(\R_src2_lo[4]~11_combout ),
	.datab(\D_iw[6]~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\E_src2[0]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[0]~16_combout ),
	.cout());
defparam \R_src2_lo[0]~16 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[0]~16 .sum_lutc_input = "datac";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\R_src2_lo[0]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

dffeas \E_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[0]~5_combout ),
	.asdata(\E_src2[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[1]~7 (
	.dataa(\E_shift_rot_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[0]~6 ),
	.combout(\E_shift_rot_cnt[1]~7_combout ),
	.cout(\E_shift_rot_cnt[1]~8 ));
defparam \E_shift_rot_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[7]~96 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(readdata_7),
	.cin(gnd),
	.combout(\F_iw[7]~96_combout ),
	.cout());
defparam \F_iw[7]~96 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~96 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~97 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_7),
	.datad(q_a_7),
	.cin(gnd),
	.combout(\F_iw[7]~97_combout ),
	.cout());
defparam \F_iw[7]~97 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~97 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~98 (
	.dataa(\F_iw[7]~96_combout ),
	.datab(\F_iw[7]~97_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_7),
	.cin(gnd),
	.combout(\F_iw[7]~98_combout ),
	.cout());
defparam \F_iw[7]~98 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~98 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~99 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[7]~98_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_71),
	.cin(gnd),
	.combout(\F_iw[7]~99_combout ),
	.cout());
defparam \F_iw[7]~99 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~99 .sum_lutc_input = "datac";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~99_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[1]~15 (
	.dataa(\R_src2_lo[4]~11_combout ),
	.datab(\D_iw[7]~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\E_src2[0]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[1]~15_combout ),
	.cout());
defparam \R_src2_lo[1]~15 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[1]~15 .sum_lutc_input = "datac";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\R_src2_lo[1]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[1]~7_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[2]~9 (
	.dataa(\E_shift_rot_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[1]~8 ),
	.combout(\E_shift_rot_cnt[2]~9_combout ),
	.cout(\E_shift_rot_cnt[2]~10 ));
defparam \E_shift_rot_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \E_shift_rot_cnt[2]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[8]~89 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_86_0),
	.datac(mem_68_0),
	.datad(readdata_8),
	.cin(gnd),
	.combout(\F_iw[8]~89_combout ),
	.cout());
defparam \F_iw[8]~89 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~90 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_8),
	.datad(q_a_8),
	.cin(gnd),
	.combout(\F_iw[8]~90_combout ),
	.cout());
defparam \F_iw[8]~90 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~91 (
	.dataa(\F_iw[8]~89_combout ),
	.datab(\F_iw[8]~90_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_8),
	.cin(gnd),
	.combout(\F_iw[8]~91_combout ),
	.cout());
defparam \F_iw[8]~91 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~92 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[8]~91_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_81),
	.cin(gnd),
	.combout(\F_iw[8]~92_combout ),
	.cout());
defparam \F_iw[8]~92 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~92 .sum_lutc_input = "datac";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~92_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[2]~14 (
	.dataa(\R_src2_lo[4]~11_combout ),
	.datab(\D_iw[8]~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datad(\E_src2[0]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[2]~14_combout ),
	.cout());
defparam \R_src2_lo[2]~14 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[2]~14 .sum_lutc_input = "datac";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\R_src2_lo[2]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[2]~9_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[3]~11 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[2]~10 ),
	.combout(\E_shift_rot_cnt[3]~11_combout ),
	.cout(\E_shift_rot_cnt[3]~12 ));
defparam \E_shift_rot_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[3]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[9]~83 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_9),
	.datad(av_readdata_pre_9),
	.cin(gnd),
	.combout(\F_iw[9]~83_combout ),
	.cout());
defparam \F_iw[9]~83 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[9]~84 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_9),
	.datad(out_data_buffer_91),
	.cin(gnd),
	.combout(\F_iw[9]~84_combout ),
	.cout());
defparam \F_iw[9]~84 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[9]~85 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[9]~83_combout ),
	.datac(\F_iw[9]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[9]~85_combout ),
	.cout());
defparam \F_iw[9]~85 .lut_mask = 16'hFEFE;
defparam \F_iw[9]~85 .sum_lutc_input = "datac";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~85_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[3]~13 (
	.dataa(\R_src2_lo[4]~11_combout ),
	.datab(\D_iw[9]~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datad(\E_src2[0]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[3]~13_combout ),
	.cout());
defparam \R_src2_lo[3]~13 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[3]~13 .sum_lutc_input = "datac";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\R_src2_lo[3]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[3]~11_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[4]~13 (
	.dataa(\E_shift_rot_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\E_shift_rot_cnt[3]~12 ),
	.combout(\E_shift_rot_cnt[4]~13_combout ),
	.cout());
defparam \E_shift_rot_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \E_shift_rot_cnt[4]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[10]~77 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_10),
	.datad(q_a_10),
	.cin(gnd),
	.combout(\F_iw[10]~77_combout ),
	.cout());
defparam \F_iw[10]~77 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~78 (
	.dataa(src_payload3),
	.datab(\F_iw[10]~77_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\F_iw[10]~78_combout ),
	.cout());
defparam \F_iw[10]~78 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~79 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[10]~78_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_101),
	.cin(gnd),
	.combout(\F_iw[10]~79_combout ),
	.cout());
defparam \F_iw[10]~79 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~79 .sum_lutc_input = "datac";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~79_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[4]~12 (
	.dataa(\R_src2_lo[4]~11_combout ),
	.datab(\D_iw[10]~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datad(\E_src2[0]~16_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~12_combout ),
	.cout());
defparam \R_src2_lo[4]~12 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[4]~12 .sum_lutc_input = "datac";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\R_src2_lo[4]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[4]~13_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cycloneive_lcell_comb \E_stall~0 (
	.dataa(\E_shift_rot_cnt[1]~q ),
	.datab(\E_shift_rot_cnt[2]~q ),
	.datac(\E_shift_rot_cnt[3]~q ),
	.datad(\E_shift_rot_cnt[4]~q ),
	.cin(gnd),
	.combout(\E_stall~0_combout ),
	.cout());
defparam \E_stall~0 .lut_mask = 16'hFFFE;
defparam \E_stall~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~1 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_shift_rot~q ),
	.datac(\E_shift_rot_cnt[0]~q ),
	.datad(\E_stall~0_combout ),
	.cin(gnd),
	.combout(\E_stall~1_combout ),
	.cout());
defparam \E_stall~1 .lut_mask = 16'hFFFE;
defparam \E_stall~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~2 (
	.dataa(\R_ctrl_ld~q ),
	.datab(\E_new_inst~q ),
	.datac(\E_valid_from_R~q ),
	.datad(\E_stall~1_combout ),
	.cin(gnd),
	.combout(\E_stall~2_combout ),
	.cout());
defparam \E_stall~2 .lut_mask = 16'hFFFE;
defparam \E_stall~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem32~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.cout());
defparam \D_ctrl_mem32~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem32~0 .sum_lutc_input = "datac";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_aligning_data_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cycloneive_lcell_comb \D_ctrl_mem16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.cout());
defparam \D_ctrl_mem16~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_mem16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[0]~0 (
	.dataa(\av_ld_align_cycle[0]~q ),
	.datab(d_read1),
	.datac(av_ld_getting_data),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~0_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[0]~0 .lut_mask = 16'h7F7F;
defparam \av_ld_align_cycle_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[0] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[1]~1 (
	.dataa(\av_ld_align_cycle[1]~q ),
	.datab(\av_ld_align_cycle[0]~q ),
	.datac(d_read1),
	.datad(av_ld_getting_data),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~1_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[1]~1 .lut_mask = 16'h6FFF;
defparam \av_ld_align_cycle_nxt[1]~1 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[1] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(\D_iw[4]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 16'h96FF;
defparam \av_ld_aligning_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(src_payload),
	.datab(d_read1),
	.datac(WideOr1),
	.datad(\av_ld_getting_data~7_combout ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 16'hFFFD;
defparam \av_ld_aligning_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~2 (
	.dataa(\D_ctrl_mem32~0_combout ),
	.datab(\av_ld_aligning_data~q ),
	.datac(\av_ld_aligning_data_nxt~0_combout ),
	.datad(\av_ld_aligning_data_nxt~1_combout ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~2_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~2 .lut_mask = 16'hF7D5;
defparam \av_ld_aligning_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~3 (
	.dataa(\E_new_inst~q ),
	.datab(\av_ld_aligning_data_nxt~2_combout ),
	.datac(\D_ctrl_mem32~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_stall~3_combout ),
	.cout());
defparam \E_stall~3 .lut_mask = 16'hEFEF;
defparam \E_stall~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~4 (
	.dataa(\av_ld_waiting_for_data_nxt~0_combout ),
	.datab(\E_stall~1_combout ),
	.datac(\E_stall~2_combout ),
	.datad(\E_stall~3_combout ),
	.cin(gnd),
	.combout(\E_stall~4_combout ),
	.cout());
defparam \E_stall~4 .lut_mask = 16'hFFFE;
defparam \E_stall~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~3 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\R_valid~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_valid_from_R~3_combout ),
	.cout());
defparam \E_valid_from_R~3 .lut_mask = 16'hFEFE;
defparam \E_valid_from_R~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~2 (
	.dataa(\E_stall~4_combout ),
	.datab(d_write1),
	.datac(av_waitrequest),
	.datad(\E_valid_from_R~3_combout ),
	.cin(gnd),
	.combout(\E_valid_from_R~2_combout ),
	.cout());
defparam \E_valid_from_R~2 .lut_mask = 16'hFFFE;
defparam \E_valid_from_R~2 .sum_lutc_input = "datac";

dffeas E_valid_from_R(
	.clk(clk_clk),
	.d(\E_valid_from_R~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cycloneive_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~0 .lut_mask = 16'h0FFF;
defparam \D_ctrl_jmp_direct~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_jmp_direct~1 (
	.dataa(\D_ctrl_jmp_direct~0_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~1_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_jmp_direct~1 .sum_lutc_input = "datac";

dffeas R_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_direct~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

dffeas R_ctrl_br(
	.clk(clk_clk),
	.d(\R_ctrl_br_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cycloneive_lcell_comb \D_ctrl_retaddr~4 (
	.dataa(\Equal62~14_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~4_combout ),
	.cout());
defparam \D_ctrl_retaddr~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_retaddr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~5 (
	.dataa(\D_ctrl_retaddr~4_combout ),
	.datab(\Equal62~8_combout ),
	.datac(\Equal62~9_combout ),
	.datad(\D_dst_regnum[4]~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~5_combout ),
	.cout());
defparam \D_ctrl_retaddr~5 .lut_mask = 16'hFEFF;
defparam \D_ctrl_retaddr~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~6 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_retaddr~5_combout ),
	.datac(\D_ctrl_force_src2_zero~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~6_combout ),
	.cout());
defparam \D_ctrl_retaddr~6 .lut_mask = 16'hF7F7;
defparam \D_ctrl_retaddr~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~9 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hFF7F;
defparam \Equal0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~7 (
	.dataa(\Equal0~13_combout ),
	.datab(\Equal0~9_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_dst_regnum[4]~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~7_combout ),
	.cout());
defparam \D_ctrl_retaddr~7 .lut_mask = 16'hFFDE;
defparam \D_ctrl_retaddr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~8 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~12_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~8_combout ),
	.cout());
defparam \D_ctrl_retaddr~8 .lut_mask = 16'hFFBE;
defparam \D_ctrl_retaddr~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~9 (
	.dataa(\Equal0~2_combout ),
	.datab(\D_ctrl_retaddr~6_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~8_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~9_combout ),
	.cout());
defparam \D_ctrl_retaddr~9 .lut_mask = 16'hBFFB;
defparam \D_ctrl_retaddr~9 .sum_lutc_input = "datac";

dffeas R_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cycloneive_lcell_comb \R_src1~11 (
	.dataa(\R_ctrl_br~q ),
	.datab(\R_valid~q ),
	.datac(\R_ctrl_retaddr~q ),
	.datad(\E_valid_from_R~q ),
	.cin(gnd),
	.combout(\R_src1~11_combout ),
	.cout());
defparam \R_src1~11 .lut_mask = 16'hFFFE;
defparam \R_src1~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[1]~12 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[1]~12_combout ),
	.cout());
defparam \R_src1[1]~12 .lut_mask = 16'hF7FF;
defparam \R_src1[1]~12 .sum_lutc_input = "datac";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\R_src1[1]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

cycloneive_lcell_comb D_op_wrctl(
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~3_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_wrctl~combout ),
	.cout());
defparam D_op_wrctl.lut_mask = 16'hFEFF;
defparam D_op_wrctl.sum_lutc_input = "datac";

dffeas R_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cycloneive_lcell_comb \W_ienable_reg_nxt~0 (
	.dataa(\D_iw[7]~q ),
	.datab(\D_iw[6]~q ),
	.datac(\R_ctrl_wrctl_inst~q ),
	.datad(\D_iw[8]~q ),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~0_combout ),
	.cout());
defparam \W_ienable_reg_nxt~0 .lut_mask = 16'hFEFF;
defparam \W_ienable_reg_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_ienable_reg_nxt~1 (
	.dataa(\E_valid_from_R~q ),
	.datab(\W_ienable_reg_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~1_combout ),
	.cout());
defparam \W_ienable_reg_nxt~1 .lut_mask = 16'hEEEE;
defparam \W_ienable_reg_nxt~1 .sum_lutc_input = "datac";

dffeas \W_ienable_reg[1] (
	.clk(clk_clk),
	.d(\E_src1[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~1_combout ),
	.q(\W_ienable_reg[1]~q ),
	.prn(vcc));
defparam \W_ienable_reg[1] .is_wysiwyg = "true";
defparam \W_ienable_reg[1] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[1]~0 (
	.dataa(\W_ienable_reg[1]~q ),
	.datab(av_readdata_9),
	.datac(av_readdata_8),
	.datad(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[1]~0_combout ),
	.cout());
defparam \W_ipending_reg_nxt[1]~0 .lut_mask = 16'hFEFF;
defparam \W_ipending_reg_nxt[1]~0 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[1] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[1]~q ),
	.prn(vcc));
defparam \W_ipending_reg[1] .is_wysiwyg = "true";
defparam \W_ipending_reg[1] .power_up = "low";

cycloneive_lcell_comb \R_src1[0]~13 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[0]~13_combout ),
	.cout());
defparam \R_src1[0]~13 .lut_mask = 16'hF7FF;
defparam \R_src1[0]~13 .sum_lutc_input = "datac";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\R_src1[0]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

dffeas \W_ienable_reg[0] (
	.clk(clk_clk),
	.d(\E_src1[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_ienable_reg_nxt~1_combout ),
	.q(\W_ienable_reg[0]~q ),
	.prn(vcc));
defparam \W_ienable_reg[0] .is_wysiwyg = "true";
defparam \W_ienable_reg[0] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[0]~1 (
	.dataa(\W_ienable_reg[0]~q ),
	.datab(dreg_1),
	.datac(gnd),
	.datad(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[0]~1_combout ),
	.cout());
defparam \W_ipending_reg_nxt[0]~1 .lut_mask = 16'hEEFF;
defparam \W_ipending_reg_nxt[0]~1 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[0] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[0]~q ),
	.prn(vcc));
defparam \W_ipending_reg[0] .is_wysiwyg = "true";
defparam \W_ipending_reg[0] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_exception~0 (
	.dataa(\Equal62~8_combout ),
	.datab(\D_op_opx_rsv63~0_combout ),
	.datac(\Equal62~9_combout ),
	.datad(\D_dst_regnum[4]~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.cout());
defparam \D_ctrl_exception~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_exception~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.cout());
defparam \D_ctrl_exception~1 .lut_mask = 16'hFBFF;
defparam \D_ctrl_exception~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~2 (
	.dataa(\D_iw[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~2_combout ),
	.cout());
defparam \D_ctrl_exception~2 .lut_mask = 16'hAAFF;
defparam \D_ctrl_exception~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~3 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_exception~0_combout ),
	.datac(\D_ctrl_exception~1_combout ),
	.datad(\D_ctrl_exception~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~3_combout ),
	.cout());
defparam \D_ctrl_exception~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~1 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~13_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~1_combout ),
	.cout());
defparam \D_dst_regnum[4]~1 .lut_mask = 16'hFEFF;
defparam \D_dst_regnum[4]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~2 (
	.dataa(\Equal0~3_combout ),
	.datab(\Equal0~2_combout ),
	.datac(\Equal0~12_combout ),
	.datad(\D_dst_regnum[4]~1_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~2_combout ),
	.cout());
defparam \D_dst_regnum[4]~2 .lut_mask = 16'hBFFF;
defparam \D_dst_regnum[4]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~4 (
	.dataa(\D_dst_regnum[4]~2_combout ),
	.datab(\D_dst_regnum[4]~3_combout ),
	.datac(\Equal0~13_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~4_combout ),
	.cout());
defparam \D_dst_regnum[4]~4 .lut_mask = 16'hEFFF;
defparam \D_dst_regnum[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~15 (
	.dataa(\D_ctrl_exception~3_combout ),
	.datab(\D_ctrl_exception~8_combout ),
	.datac(\D_ctrl_exception~14_combout ),
	.datad(\D_dst_regnum[4]~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~15_combout ),
	.cout());
defparam \D_ctrl_exception~15 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~15 .sum_lutc_input = "datac";

dffeas R_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cycloneive_lcell_comb \D_ctrl_break~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\D_iw[16]~q ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.cout());
defparam \D_ctrl_break~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_break~0 .sum_lutc_input = "datac";

dffeas R_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

cycloneive_lcell_comb \F_pc_no_crst_nxt[25]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\R_ctrl_exception~q ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[25]~5_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[25]~5 .lut_mask = 16'h0FFF;
defparam \F_pc_no_crst_nxt[25]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal132~2 (
	.dataa(\D_iw[6]~q ),
	.datab(\R_ctrl_wrctl_inst~q ),
	.datac(\D_iw[8]~q ),
	.datad(\D_iw[7]~q ),
	.cin(gnd),
	.combout(\Equal132~2_combout ),
	.cout());
defparam \Equal132~2 .lut_mask = 16'hEFFF;
defparam \Equal132~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_estatus_reg~q ),
	.datac(\Equal132~2_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 16'hACFF;
defparam \W_estatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~1 (
	.dataa(\W_estatus_reg_inst_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\W_status_reg_pie~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~1 .lut_mask = 16'hFEFE;
defparam \W_estatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_estatus_reg(
	.clk(clk_clk),
	.d(\W_estatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

cycloneive_lcell_comb \Equal132~1 (
	.dataa(\D_iw[7]~q ),
	.datab(\R_ctrl_wrctl_inst~q ),
	.datac(\D_iw[8]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\Equal132~1_combout ),
	.cout());
defparam \Equal132~1 .lut_mask = 16'hEFFF;
defparam \Equal132~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_bstatus_reg~q ),
	.datac(\Equal132~1_combout ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 16'hACFF;
defparam \W_bstatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~1 (
	.dataa(\W_bstatus_reg_inst_nxt~0_combout ),
	.datab(\R_ctrl_break~q ),
	.datac(\W_status_reg_pie~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~1 .lut_mask = 16'hFEFE;
defparam \W_bstatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

dffeas W_bstatus_reg(
	.clk(clk_clk),
	.d(\W_bstatus_reg_inst_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cycloneive_lcell_comb \Equal132~0 (
	.dataa(\R_ctrl_wrctl_inst~q ),
	.datab(\D_iw[8]~q ),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\Equal132~0_combout ),
	.cout());
defparam \Equal132~0 .lut_mask = 16'hBFFF;
defparam \Equal132~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_status_reg_pie~q ),
	.datac(gnd),
	.datad(\Equal132~0_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 16'hAACC;
defparam \W_status_reg_pie_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~0_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\Equal62~10_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_op_eret(
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~10_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_eret~combout ),
	.cout());
defparam D_op_eret.lut_mask = 16'hEFFF;
defparam D_op_eret.sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\W_estatus_reg~q ),
	.datac(\W_status_reg_pie_inst_nxt~1_combout ),
	.datad(\D_op_eret~combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 16'hFAFC;
defparam \W_status_reg_pie_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cycloneive_lcell_comb \D_iw[26]~0 (
	.dataa(gnd),
	.datab(\W_ipending_reg[1]~q ),
	.datac(\W_ipending_reg[0]~q ),
	.datad(\W_status_reg_pie~q ),
	.cin(gnd),
	.combout(\D_iw[26]~0_combout ),
	.cout());
defparam \D_iw[26]~0 .lut_mask = 16'h3FFF;
defparam \D_iw[26]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_iw[26]~1 (
	.dataa(\D_iw[26]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(gnd),
	.datad(\hbreak_req~0_combout ),
	.cin(gnd),
	.combout(\D_iw[26]~1_combout ),
	.cout());
defparam \D_iw[26]~1 .lut_mask = 16'hEEFF;
defparam \D_iw[26]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[11]~25 (
	.dataa(src1_valid1),
	.datab(av_readdata_pre_111),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[11]~25_combout ),
	.cout());
defparam \F_iw[11]~25 .lut_mask = 16'hEEFF;
defparam \F_iw[11]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[11]~26 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_111),
	.datad(out_data_buffer_112),
	.cin(gnd),
	.combout(\F_iw[11]~26_combout ),
	.cout());
defparam \F_iw[11]~26 .lut_mask = 16'hFFFE;
defparam \F_iw[11]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[11]~27 (
	.dataa(\F_iw[11]~25_combout ),
	.datab(\F_iw[11]~26_combout ),
	.datac(src1_valid2),
	.datad(q_a_11),
	.cin(gnd),
	.combout(\F_iw[11]~27_combout ),
	.cout());
defparam \F_iw[11]~27 .lut_mask = 16'hFFFE;
defparam \F_iw[11]~27 .sum_lutc_input = "datac";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cycloneive_lcell_comb \Equal62~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~0_combout ),
	.cout());
defparam \Equal62~0 .lut_mask = 16'h7FFF;
defparam \Equal62~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hFFBF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~8 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~5_combout ),
	.datad(\D_ctrl_alu_force_xor~14_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~8_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~8 .lut_mask = 16'h27FF;
defparam \D_ctrl_alu_subtract~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~9 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_alu_subtract~8_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~9_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~9 .lut_mask = 16'hEEFF;
defparam \D_ctrl_alu_subtract~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~5 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~5_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~5 .lut_mask = 16'hFF96;
defparam \D_ctrl_alu_subtract~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~10 (
	.dataa(\D_ctrl_alu_subtract~5_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~10_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~10 .lut_mask = 16'hBFBF;
defparam \D_ctrl_alu_subtract~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_alu_sub~0 (
	.dataa(\R_valid~q ),
	.datab(\D_ctrl_alu_subtract~9_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_subtract~10_combout ),
	.cin(gnd),
	.combout(\E_alu_sub~0_combout ),
	.cout());
defparam \E_alu_sub~0 .lut_mask = 16'hFFFE;
defparam \E_alu_sub~0 .sum_lutc_input = "datac";

dffeas E_alu_sub(
	.clk(clk_clk),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cycloneive_lcell_comb \F_iw[21]~46 (
	.dataa(src1_valid1),
	.datab(av_readdata_pre_21),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[21]~46_combout ),
	.cout());
defparam \F_iw[21]~46 .lut_mask = 16'hEEFF;
defparam \F_iw[21]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[21]~47 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_211),
	.datad(out_data_buffer_212),
	.cin(gnd),
	.combout(\F_iw[21]~47_combout ),
	.cout());
defparam \F_iw[21]~47 .lut_mask = 16'hFFFE;
defparam \F_iw[21]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[21]~48 (
	.dataa(\F_iw[21]~46_combout ),
	.datab(\F_iw[21]~47_combout ),
	.datac(src1_valid2),
	.datad(q_a_21),
	.cin(gnd),
	.combout(\F_iw[21]~48_combout ),
	.cout());
defparam \F_iw[21]~48 .lut_mask = 16'hFFFE;
defparam \F_iw[21]~48 .sum_lutc_input = "datac";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cycloneive_lcell_comb \E_src2[28]~0 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[28]~0_combout ),
	.cout());
defparam \E_src2[28]~0 .lut_mask = 16'hAACC;
defparam \E_src2[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~49 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_18),
	.datad(q_a_18),
	.cin(gnd),
	.combout(\F_iw[18]~49_combout ),
	.cout());
defparam \F_iw[18]~49 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~50 (
	.dataa(src_payload3),
	.datab(\F_iw[18]~49_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_18),
	.cin(gnd),
	.combout(\F_iw[18]~50_combout ),
	.cout());
defparam \F_iw[18]~50 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~51 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[18]~50_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_181),
	.cin(gnd),
	.combout(\F_iw[18]~51_combout ),
	.cout());
defparam \F_iw[18]~51 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~52 (
	.dataa(\F_iw[18]~51_combout ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\F_iw[18]~52_combout ),
	.cout());
defparam \F_iw[18]~52 .lut_mask = 16'hEEFF;
defparam \F_iw[18]~52 .sum_lutc_input = "datac";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hF7FF;
defparam \Equal0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~6_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~3 .lut_mask = 16'hFAFC;
defparam \D_ctrl_unsigned_lo_imm16~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~10 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
defparam \Equal0~10 .lut_mask = 16'hFFF7;
defparam \Equal0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_logic~0 (
	.dataa(gnd),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~9_combout ),
	.datad(\Equal0~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.cout());
defparam \D_ctrl_logic~0 .lut_mask = 16'h3FFF;
defparam \D_ctrl_logic~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~4 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_unsigned_lo_imm16~4 .sum_lutc_input = "datac";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cycloneive_lcell_comb \R_src2_hi~0 (
	.dataa(\R_ctrl_force_src2_zero~q ),
	.datab(\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_hi~0_combout ),
	.cout());
defparam \R_src2_hi~0 .lut_mask = 16'hEEEE;
defparam \R_src2_hi~0 .sum_lutc_input = "datac";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\E_src2[28]~0_combout ),
	.asdata(\D_iw[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[28]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_valid_from_R~q ),
	.datad(\R_ctrl_jmp_direct~q ),
	.cin(gnd),
	.combout(\R_src1~10_combout ),
	.cout());
defparam \R_src1~10 .lut_mask = 16'h0FFF;
defparam \R_src1~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[28]~0 (
	.dataa(F_pc_26),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[28]~0_combout ),
	.cout());
defparam \E_src1[28]~0 .lut_mask = 16'hCC55;
defparam \E_src1[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[0]~0 (
	.dataa(F_pc_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\F_pc_plus_one[0]~0_combout ),
	.cout(\F_pc_plus_one[0]~1 ));
defparam \F_pc_plus_one[0]~0 .lut_mask = 16'h55AA;
defparam \F_pc_plus_one[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[1]~2 (
	.dataa(F_pc_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[0]~1 ),
	.combout(\F_pc_plus_one[1]~2_combout ),
	.cout(\F_pc_plus_one[1]~3 ));
defparam \F_pc_plus_one[1]~2 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[2]~4 (
	.dataa(F_pc_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[1]~3 ),
	.combout(\F_pc_plus_one[2]~4_combout ),
	.cout(\F_pc_plus_one[2]~5 ));
defparam \F_pc_plus_one[2]~4 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[3]~6 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[2]~5 ),
	.combout(\F_pc_plus_one[3]~6_combout ),
	.cout(\F_pc_plus_one[3]~7 ));
defparam \F_pc_plus_one[3]~6 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[4]~8 (
	.dataa(F_pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[3]~7 ),
	.combout(\F_pc_plus_one[4]~8_combout ),
	.cout(\F_pc_plus_one[4]~9 ));
defparam \F_pc_plus_one[4]~8 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[4]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[5]~10 (
	.dataa(F_pc_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[4]~9 ),
	.combout(\F_pc_plus_one[5]~10_combout ),
	.cout(\F_pc_plus_one[5]~11 ));
defparam \F_pc_plus_one[5]~10 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[6]~12 (
	.dataa(F_pc_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[5]~11 ),
	.combout(\F_pc_plus_one[6]~12_combout ),
	.cout(\F_pc_plus_one[6]~13 ));
defparam \F_pc_plus_one[6]~12 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[7]~14 (
	.dataa(F_pc_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[6]~13 ),
	.combout(\F_pc_plus_one[7]~14_combout ),
	.cout(\F_pc_plus_one[7]~15 ));
defparam \F_pc_plus_one[7]~14 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[8]~16 (
	.dataa(F_pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[7]~15 ),
	.combout(\F_pc_plus_one[8]~16_combout ),
	.cout(\F_pc_plus_one[8]~17 ));
defparam \F_pc_plus_one[8]~16 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[9]~18 (
	.dataa(F_pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[8]~17 ),
	.combout(\F_pc_plus_one[9]~18_combout ),
	.cout(\F_pc_plus_one[9]~19 ));
defparam \F_pc_plus_one[9]~18 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[9]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[10]~20 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[9]~19 ),
	.combout(\F_pc_plus_one[10]~20_combout ),
	.cout(\F_pc_plus_one[10]~21 ));
defparam \F_pc_plus_one[10]~20 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[10]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[11]~22 (
	.dataa(F_pc_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[10]~21 ),
	.combout(\F_pc_plus_one[11]~22_combout ),
	.cout(\F_pc_plus_one[11]~23 ));
defparam \F_pc_plus_one[11]~22 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[11]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[12]~24 (
	.dataa(F_pc_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[11]~23 ),
	.combout(\F_pc_plus_one[12]~24_combout ),
	.cout(\F_pc_plus_one[12]~25 ));
defparam \F_pc_plus_one[12]~24 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[12]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[13]~26 (
	.dataa(F_pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[12]~25 ),
	.combout(\F_pc_plus_one[13]~26_combout ),
	.cout(\F_pc_plus_one[13]~27 ));
defparam \F_pc_plus_one[13]~26 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[13]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[14]~28 (
	.dataa(F_pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[13]~27 ),
	.combout(\F_pc_plus_one[14]~28_combout ),
	.cout(\F_pc_plus_one[14]~29 ));
defparam \F_pc_plus_one[14]~28 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[14]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[15]~30 (
	.dataa(F_pc_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[14]~29 ),
	.combout(\F_pc_plus_one[15]~30_combout ),
	.cout(\F_pc_plus_one[15]~31 ));
defparam \F_pc_plus_one[15]~30 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[15]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[16]~32 (
	.dataa(F_pc_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[15]~31 ),
	.combout(\F_pc_plus_one[16]~32_combout ),
	.cout(\F_pc_plus_one[16]~33 ));
defparam \F_pc_plus_one[16]~32 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[16]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[17]~34 (
	.dataa(F_pc_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[16]~33 ),
	.combout(\F_pc_plus_one[17]~34_combout ),
	.cout(\F_pc_plus_one[17]~35 ));
defparam \F_pc_plus_one[17]~34 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[17]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[18]~36 (
	.dataa(F_pc_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[17]~35 ),
	.combout(\F_pc_plus_one[18]~36_combout ),
	.cout(\F_pc_plus_one[18]~37 ));
defparam \F_pc_plus_one[18]~36 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[18]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[19]~38 (
	.dataa(F_pc_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[18]~37 ),
	.combout(\F_pc_plus_one[19]~38_combout ),
	.cout(\F_pc_plus_one[19]~39 ));
defparam \F_pc_plus_one[19]~38 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[19]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[20]~40 (
	.dataa(F_pc_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[19]~39 ),
	.combout(\F_pc_plus_one[20]~40_combout ),
	.cout(\F_pc_plus_one[20]~41 ));
defparam \F_pc_plus_one[20]~40 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[20]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[21]~42 (
	.dataa(F_pc_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[20]~41 ),
	.combout(\F_pc_plus_one[21]~42_combout ),
	.cout(\F_pc_plus_one[21]~43 ));
defparam \F_pc_plus_one[21]~42 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[21]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[22]~44 (
	.dataa(F_pc_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[21]~43 ),
	.combout(\F_pc_plus_one[22]~44_combout ),
	.cout(\F_pc_plus_one[22]~45 ));
defparam \F_pc_plus_one[22]~44 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[22]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[23]~46 (
	.dataa(F_pc_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[22]~45 ),
	.combout(\F_pc_plus_one[23]~46_combout ),
	.cout(\F_pc_plus_one[23]~47 ));
defparam \F_pc_plus_one[23]~46 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[23]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[24]~48 (
	.dataa(F_pc_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[23]~47 ),
	.combout(\F_pc_plus_one[24]~48_combout ),
	.cout(\F_pc_plus_one[24]~49 ));
defparam \F_pc_plus_one[24]~48 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[24]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[25]~50 (
	.dataa(F_pc_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[24]~49 ),
	.combout(\F_pc_plus_one[25]~50_combout ),
	.cout(\F_pc_plus_one[25]~51 ));
defparam \F_pc_plus_one[25]~50 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[25]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[26]~52 (
	.dataa(F_pc_26),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\F_pc_plus_one[25]~51 ),
	.combout(\F_pc_plus_one[26]~52_combout ),
	.cout());
defparam \F_pc_plus_one[26]~52 .lut_mask = 16'h5A5A;
defparam \F_pc_plus_one[26]~52 .sum_lutc_input = "cin";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\E_src1[28]~0_combout ),
	.asdata(\F_pc_plus_one[26]~52_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

cycloneive_lcell_comb \E_src2[27]~1 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[27]~1_combout ),
	.cout());
defparam \E_src2[27]~1 .lut_mask = 16'hAACC;
defparam \E_src2[27]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~53 (
	.dataa(src1_valid),
	.datab(src1_valid1),
	.datac(av_readdata_pre_17),
	.datad(readdata_17),
	.cin(gnd),
	.combout(\F_iw[17]~53_combout ),
	.cout());
defparam \F_iw[17]~53 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~54 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_17),
	.datad(q_a_17),
	.cin(gnd),
	.combout(\F_iw[17]~54_combout ),
	.cout());
defparam \F_iw[17]~54 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~55 (
	.dataa(\F_iw[17]~53_combout ),
	.datab(\F_iw[17]~54_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_171),
	.cin(gnd),
	.combout(\F_iw[17]~55_combout ),
	.cout());
defparam \F_iw[17]~55 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~111 (
	.dataa(\D_iw[26]~0_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\F_iw[17]~55_combout ),
	.cin(gnd),
	.combout(\F_iw[17]~111_combout ),
	.cout());
defparam \F_iw[17]~111 .lut_mask = 16'hFFDF;
defparam \F_iw[17]~111 .sum_lutc_input = "datac";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~111_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\E_src2[27]~1_combout ),
	.asdata(\D_iw[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[27]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~56 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_31),
	.datad(av_readdata_pre_31),
	.cin(gnd),
	.combout(\F_iw[31]~56_combout ),
	.cout());
defparam \F_iw[31]~56 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~57 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_311),
	.datad(out_data_buffer_312),
	.cin(gnd),
	.combout(\F_iw[31]~57_combout ),
	.cout());
defparam \F_iw[31]~57 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~58 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[31]~56_combout ),
	.datac(\F_iw[31]~57_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[31]~58_combout ),
	.cout());
defparam \F_iw[31]~58 .lut_mask = 16'hFEFE;
defparam \F_iw[31]~58 .sum_lutc_input = "datac";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~58_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cycloneive_lcell_comb \E_src1[27]~1 (
	.dataa(\D_iw[31]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[27]~1_combout ),
	.cout());
defparam \E_src1[27]~1 .lut_mask = 16'hAACC;
defparam \E_src1[27]~1 .sum_lutc_input = "datac";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\E_src1[27]~1_combout ),
	.asdata(\F_pc_plus_one[25]~50_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

cycloneive_lcell_comb \E_src2[26]~2 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[26]~2_combout ),
	.cout());
defparam \E_src2[26]~2 .lut_mask = 16'hAACC;
defparam \E_src2[26]~2 .sum_lutc_input = "datac";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\E_src2[26]~2_combout ),
	.asdata(\D_iw[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[26]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~59 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_30),
	.datad(q_a_30),
	.cin(gnd),
	.combout(\F_iw[30]~59_combout ),
	.cout());
defparam \F_iw[30]~59 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~60 (
	.dataa(src_payload3),
	.datab(\F_iw[30]~59_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\F_iw[30]~60_combout ),
	.cout());
defparam \F_iw[30]~60 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~61 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[30]~60_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_301),
	.cin(gnd),
	.combout(\F_iw[30]~61_combout ),
	.cout());
defparam \F_iw[30]~61 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~61 .sum_lutc_input = "datac";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~61_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

cycloneive_lcell_comb \E_src1[26]~2 (
	.dataa(\D_iw[30]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[26]~2_combout ),
	.cout());
defparam \E_src1[26]~2 .lut_mask = 16'hAACC;
defparam \E_src1[26]~2 .sum_lutc_input = "datac";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\E_src1[26]~2_combout ),
	.asdata(\F_pc_plus_one[24]~48_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

cycloneive_lcell_comb \E_src2[25]~3 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[25]~3_combout ),
	.cout());
defparam \E_src2[25]~3 .lut_mask = 16'hAACC;
defparam \E_src2[25]~3 .sum_lutc_input = "datac";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\E_src2[25]~3_combout ),
	.asdata(\D_iw[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cycloneive_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[25]~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~62 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_29),
	.datad(av_readdata_pre_29),
	.cin(gnd),
	.combout(\F_iw[29]~62_combout ),
	.cout());
defparam \F_iw[29]~62 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~63 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_29),
	.datad(out_data_buffer_291),
	.cin(gnd),
	.combout(\F_iw[29]~63_combout ),
	.cout());
defparam \F_iw[29]~63 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~64 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[29]~62_combout ),
	.datac(\F_iw[29]~63_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[29]~64_combout ),
	.cout());
defparam \F_iw[29]~64 .lut_mask = 16'hFEFE;
defparam \F_iw[29]~64 .sum_lutc_input = "datac";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

cycloneive_lcell_comb \E_src1[25]~3 (
	.dataa(\D_iw[29]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[25]~3_combout ),
	.cout());
defparam \E_src1[25]~3 .lut_mask = 16'hAACC;
defparam \E_src1[25]~3 .sum_lutc_input = "datac";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\E_src1[25]~3_combout ),
	.asdata(\F_pc_plus_one[23]~46_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

cycloneive_lcell_comb \E_src2[24]~4 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[24]~4_combout ),
	.cout());
defparam \E_src2[24]~4 .lut_mask = 16'hAACC;
defparam \E_src2[24]~4 .sum_lutc_input = "datac";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\E_src2[24]~4_combout ),
	.asdata(\D_iw[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[24]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~65 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_28),
	.datad(q_a_28),
	.cin(gnd),
	.combout(\F_iw[28]~65_combout ),
	.cout());
defparam \F_iw[28]~65 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~66 (
	.dataa(src_payload3),
	.datab(\F_iw[28]~65_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\F_iw[28]~66_combout ),
	.cout());
defparam \F_iw[28]~66 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~67 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[28]~66_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_281),
	.cin(gnd),
	.combout(\F_iw[28]~67_combout ),
	.cout());
defparam \F_iw[28]~67 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~67 .sum_lutc_input = "datac";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~67_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

cycloneive_lcell_comb \E_src1[24]~4 (
	.dataa(\D_iw[28]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[24]~4_combout ),
	.cout());
defparam \E_src1[24]~4 .lut_mask = 16'hAACC;
defparam \E_src1[24]~4 .sum_lutc_input = "datac";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\E_src1[24]~4_combout ),
	.asdata(\F_pc_plus_one[22]~44_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

cycloneive_lcell_comb \E_src2[23]~5 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[23]~5_combout ),
	.cout());
defparam \E_src2[23]~5 .lut_mask = 16'hAACC;
defparam \E_src2[23]~5 .sum_lutc_input = "datac";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\E_src2[23]~5_combout ),
	.asdata(\D_iw[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cycloneive_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[23]~q ),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~68 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_27),
	.datad(av_readdata_pre_27),
	.cin(gnd),
	.combout(\F_iw[27]~68_combout ),
	.cout());
defparam \F_iw[27]~68 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~69 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_27),
	.datad(out_data_buffer_271),
	.cin(gnd),
	.combout(\F_iw[27]~69_combout ),
	.cout());
defparam \F_iw[27]~69 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~70 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[27]~68_combout ),
	.datac(\F_iw[27]~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[27]~70_combout ),
	.cout());
defparam \F_iw[27]~70 .lut_mask = 16'hFEFE;
defparam \F_iw[27]~70 .sum_lutc_input = "datac";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~70_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cycloneive_lcell_comb \E_src1[23]~5 (
	.dataa(\D_iw[27]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[23]~5_combout ),
	.cout());
defparam \E_src1[23]~5 .lut_mask = 16'hAACC;
defparam \E_src1[23]~5 .sum_lutc_input = "datac";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\E_src1[23]~5_combout ),
	.asdata(\F_pc_plus_one[21]~42_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

cycloneive_lcell_comb \E_src2[22]~6 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[22]~6_combout ),
	.cout());
defparam \E_src2[22]~6 .lut_mask = 16'hAACC;
defparam \E_src2[22]~6 .sum_lutc_input = "datac";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\E_src2[22]~6_combout ),
	.asdata(\D_iw[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[22]~q ),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~71 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_26),
	.datad(q_a_26),
	.cin(gnd),
	.combout(\F_iw[26]~71_combout ),
	.cout());
defparam \F_iw[26]~71 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~72 (
	.dataa(src_payload3),
	.datab(\F_iw[26]~71_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\F_iw[26]~72_combout ),
	.cout());
defparam \F_iw[26]~72 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~73 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[26]~72_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_261),
	.cin(gnd),
	.combout(\F_iw[26]~73_combout ),
	.cout());
defparam \F_iw[26]~73 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~73 .sum_lutc_input = "datac";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~73_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cycloneive_lcell_comb \E_src1[22]~6 (
	.dataa(\D_iw[26]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[22]~6_combout ),
	.cout());
defparam \E_src1[22]~6 .lut_mask = 16'hAACC;
defparam \E_src1[22]~6 .sum_lutc_input = "datac";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\E_src1[22]~6_combout ),
	.asdata(\F_pc_plus_one[20]~40_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

cycloneive_lcell_comb \E_src2[21]~7 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[21]~7_combout ),
	.cout());
defparam \E_src2[21]~7 .lut_mask = 16'hAACC;
defparam \E_src2[21]~7 .sum_lutc_input = "datac";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\E_src2[21]~7_combout ),
	.asdata(\D_iw[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cycloneive_lcell_comb \Add1~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[21]~q ),
	.cin(gnd),
	.combout(\Add1~7_combout ),
	.cout());
defparam \Add1~7 .lut_mask = 16'h0FF0;
defparam \Add1~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~74 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_25),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\F_iw[25]~74_combout ),
	.cout());
defparam \F_iw[25]~74 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~75 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_25),
	.datad(out_data_buffer_251),
	.cin(gnd),
	.combout(\F_iw[25]~75_combout ),
	.cout());
defparam \F_iw[25]~75 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~76 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[25]~74_combout ),
	.datac(\F_iw[25]~75_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[25]~76_combout ),
	.cout());
defparam \F_iw[25]~76 .lut_mask = 16'hFEFE;
defparam \F_iw[25]~76 .sum_lutc_input = "datac";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~76_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cycloneive_lcell_comb \E_src1[21]~7 (
	.dataa(\D_iw[25]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[21]~7_combout ),
	.cout());
defparam \E_src1[21]~7 .lut_mask = 16'hAACC;
defparam \E_src1[21]~7 .sum_lutc_input = "datac";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\E_src1[21]~7_combout ),
	.asdata(\F_pc_plus_one[19]~38_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

cycloneive_lcell_comb \E_src2[20]~8 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[20]~8_combout ),
	.cout());
defparam \E_src2[20]~8 .lut_mask = 16'hAACC;
defparam \E_src2[20]~8 .sum_lutc_input = "datac";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\E_src2[20]~8_combout ),
	.asdata(\D_iw[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[20]~q ),
	.cin(gnd),
	.combout(\Add1~8_combout ),
	.cout());
defparam \Add1~8 .lut_mask = 16'h0FF0;
defparam \Add1~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~80 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_24),
	.datad(q_a_24),
	.cin(gnd),
	.combout(\F_iw[24]~80_combout ),
	.cout());
defparam \F_iw[24]~80 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~81 (
	.dataa(src_payload3),
	.datab(\F_iw[24]~80_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\F_iw[24]~81_combout ),
	.cout());
defparam \F_iw[24]~81 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~82 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[24]~81_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_241),
	.cin(gnd),
	.combout(\F_iw[24]~82_combout ),
	.cout());
defparam \F_iw[24]~82 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~82 .sum_lutc_input = "datac";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~82_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cycloneive_lcell_comb \E_src1[20]~8 (
	.dataa(\D_iw[24]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[20]~8_combout ),
	.cout());
defparam \E_src1[20]~8 .lut_mask = 16'hAACC;
defparam \E_src1[20]~8 .sum_lutc_input = "datac";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\E_src1[20]~8_combout ),
	.asdata(\F_pc_plus_one[18]~36_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

cycloneive_lcell_comb \E_src2[19]~9 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[19]~9_combout ),
	.cout());
defparam \E_src2[19]~9 .lut_mask = 16'hAACC;
defparam \E_src2[19]~9 .sum_lutc_input = "datac";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\E_src2[19]~9_combout ),
	.asdata(\D_iw[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cycloneive_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[19]~q ),
	.cin(gnd),
	.combout(\Add1~9_combout ),
	.cout());
defparam \Add1~9 .lut_mask = 16'h0FF0;
defparam \Add1~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~86 (
	.dataa(src1_valid1),
	.datab(src1_valid2),
	.datac(q_a_23),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\F_iw[23]~86_combout ),
	.cout());
defparam \F_iw[23]~86 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~87 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_23),
	.datad(out_data_buffer_231),
	.cin(gnd),
	.combout(\F_iw[23]~87_combout ),
	.cout());
defparam \F_iw[23]~87 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~87 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~88 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[23]~86_combout ),
	.datac(\F_iw[23]~87_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_iw[23]~88_combout ),
	.cout());
defparam \F_iw[23]~88 .lut_mask = 16'hFEFE;
defparam \F_iw[23]~88 .sum_lutc_input = "datac";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~88_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cycloneive_lcell_comb \E_src1[19]~9 (
	.dataa(\D_iw[23]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[19]~9_combout ),
	.cout());
defparam \E_src1[19]~9 .lut_mask = 16'hAACC;
defparam \E_src1[19]~9 .sum_lutc_input = "datac";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\E_src1[19]~9_combout ),
	.asdata(\F_pc_plus_one[17]~34_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

cycloneive_lcell_comb \E_src2[18]~10 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[18]~10_combout ),
	.cout());
defparam \E_src2[18]~10 .lut_mask = 16'hAACC;
defparam \E_src2[18]~10 .sum_lutc_input = "datac";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\E_src2[18]~10_combout ),
	.asdata(\D_iw[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cycloneive_lcell_comb \Add1~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[18]~q ),
	.cin(gnd),
	.combout(\Add1~10_combout ),
	.cout());
defparam \Add1~10 .lut_mask = 16'h0FF0;
defparam \Add1~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~93 (
	.dataa(src1_valid2),
	.datab(out_valid2),
	.datac(out_data_buffer_22),
	.datad(q_a_22),
	.cin(gnd),
	.combout(\F_iw[22]~93_combout ),
	.cout());
defparam \F_iw[22]~93 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~93 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~94 (
	.dataa(src_payload3),
	.datab(\F_iw[22]~93_combout ),
	.datac(src1_valid1),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\F_iw[22]~94_combout ),
	.cout());
defparam \F_iw[22]~94 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~94 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~95 (
	.dataa(\D_iw[26]~1_combout ),
	.datab(\F_iw[22]~94_combout ),
	.datac(out_valid3),
	.datad(out_data_buffer_221),
	.cin(gnd),
	.combout(\F_iw[22]~95_combout ),
	.cout());
defparam \F_iw[22]~95 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~95 .sum_lutc_input = "datac";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~95_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cycloneive_lcell_comb \E_src1[18]~10 (
	.dataa(\D_iw[22]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[18]~10_combout ),
	.cout());
defparam \E_src1[18]~10 .lut_mask = 16'hAACC;
defparam \E_src1[18]~10 .sum_lutc_input = "datac";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\E_src1[18]~10_combout ),
	.asdata(\F_pc_plus_one[16]~32_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

cycloneive_lcell_comb \E_src2[17]~11 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[17]~11_combout ),
	.cout());
defparam \E_src2[17]~11 .lut_mask = 16'hAACC;
defparam \E_src2[17]~11 .sum_lutc_input = "datac";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\E_src2[17]~11_combout ),
	.asdata(\D_iw[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cycloneive_lcell_comb \Add1~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[17]~q ),
	.cin(gnd),
	.combout(\Add1~11_combout ),
	.cout());
defparam \Add1~11 .lut_mask = 16'h0FF0;
defparam \Add1~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[17]~11 (
	.dataa(\D_iw[21]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[17]~11_combout ),
	.cout());
defparam \E_src1[17]~11 .lut_mask = 16'hAACC;
defparam \E_src1[17]~11 .sum_lutc_input = "datac";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\E_src1[17]~11_combout ),
	.asdata(\F_pc_plus_one[15]~30_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

cycloneive_lcell_comb \E_src2[16]~12 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[16]~12_combout ),
	.cout());
defparam \E_src2[16]~12 .lut_mask = 16'hAACC;
defparam \E_src2[16]~12 .sum_lutc_input = "datac";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\E_src2[16]~12_combout ),
	.asdata(\D_iw[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cycloneive_lcell_comb \Add1~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[16]~q ),
	.cin(gnd),
	.combout(\Add1~12_combout ),
	.cout());
defparam \Add1~12 .lut_mask = 16'h0FF0;
defparam \Add1~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~104 (
	.dataa(src1_valid1),
	.datab(av_readdata_pre_20),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[20]~104_combout ),
	.cout());
defparam \F_iw[20]~104 .lut_mask = 16'hEEFF;
defparam \F_iw[20]~104 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~105 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_20),
	.datad(out_data_buffer_201),
	.cin(gnd),
	.combout(\F_iw[20]~105_combout ),
	.cout());
defparam \F_iw[20]~105 .lut_mask = 16'hFFFE;
defparam \F_iw[20]~105 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~106 (
	.dataa(\F_iw[20]~104_combout ),
	.datab(\F_iw[20]~105_combout ),
	.datac(src1_valid2),
	.datad(q_a_20),
	.cin(gnd),
	.combout(\F_iw[20]~106_combout ),
	.cout());
defparam \F_iw[20]~106 .lut_mask = 16'hFFFE;
defparam \F_iw[20]~106 .sum_lutc_input = "datac";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~106_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cycloneive_lcell_comb \E_src1[16]~12 (
	.dataa(\D_iw[20]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[16]~12_combout ),
	.cout());
defparam \E_src1[16]~12 .lut_mask = 16'hAACC;
defparam \E_src1[16]~12 .sum_lutc_input = "datac";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\E_src1[16]~12_combout ),
	.asdata(\F_pc_plus_one[14]~28_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

cycloneive_lcell_comb \E_src2[5]~15 (
	.dataa(\R_ctrl_src_imm5_shift_rot~q ),
	.datab(\R_ctrl_hi_imm16~q ),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[5]~15_combout ),
	.cout());
defparam \E_src2[5]~15 .lut_mask = 16'hFEFE;
defparam \E_src2[5]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[15]~0 (
	.dataa(\D_iw[21]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[15]~0_combout ),
	.cout());
defparam \R_src2_lo[15]~0 .lut_mask = 16'hACFF;
defparam \R_src2_lo[15]~0 .sum_lutc_input = "datac";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\R_src2_lo[15]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cycloneive_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[15]~q ),
	.cin(gnd),
	.combout(\Add1~13_combout ),
	.cout());
defparam \Add1~13 .lut_mask = 16'h0FF0;
defparam \Add1~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~107 (
	.dataa(src1_valid1),
	.datab(av_readdata_pre_19),
	.datac(gnd),
	.datad(\D_iw[26]~1_combout ),
	.cin(gnd),
	.combout(\F_iw[19]~107_combout ),
	.cout());
defparam \F_iw[19]~107 .lut_mask = 16'hEEFF;
defparam \F_iw[19]~107 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~108 (
	.dataa(out_valid2),
	.datab(out_valid3),
	.datac(out_data_buffer_19),
	.datad(out_data_buffer_191),
	.cin(gnd),
	.combout(\F_iw[19]~108_combout ),
	.cout());
defparam \F_iw[19]~108 .lut_mask = 16'hFFFE;
defparam \F_iw[19]~108 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~109 (
	.dataa(\F_iw[19]~107_combout ),
	.datab(\F_iw[19]~108_combout ),
	.datac(src1_valid2),
	.datad(q_a_19),
	.cin(gnd),
	.combout(\F_iw[19]~109_combout ),
	.cout());
defparam \F_iw[19]~109 .lut_mask = 16'hFFFE;
defparam \F_iw[19]~109 .sum_lutc_input = "datac";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~109_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cycloneive_lcell_comb \E_src1[15]~13 (
	.dataa(\D_iw[19]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[15]~13_combout ),
	.cout());
defparam \E_src1[15]~13 .lut_mask = 16'hAACC;
defparam \E_src1[15]~13 .sum_lutc_input = "datac";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\E_src1[15]~13_combout ),
	.asdata(\F_pc_plus_one[13]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[14]~1 (
	.dataa(\D_iw[20]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[14]~1_combout ),
	.cout());
defparam \R_src2_lo[14]~1 .lut_mask = 16'hACFF;
defparam \R_src2_lo[14]~1 .sum_lutc_input = "datac";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\R_src2_lo[14]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cycloneive_lcell_comb \Add1~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[14]~q ),
	.cin(gnd),
	.combout(\Add1~14_combout ),
	.cout());
defparam \Add1~14 .lut_mask = 16'h0FF0;
defparam \Add1~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[14]~14 (
	.dataa(\D_iw[18]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[14]~14_combout ),
	.cout());
defparam \E_src1[14]~14 .lut_mask = 16'hAACC;
defparam \E_src1[14]~14 .sum_lutc_input = "datac";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\E_src1[14]~14_combout ),
	.asdata(\F_pc_plus_one[12]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[13]~2 (
	.dataa(\D_iw[19]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[13]~2_combout ),
	.cout());
defparam \R_src2_lo[13]~2 .lut_mask = 16'hACFF;
defparam \R_src2_lo[13]~2 .sum_lutc_input = "datac";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\R_src2_lo[13]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cycloneive_lcell_comb \Add1~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[13]~q ),
	.cin(gnd),
	.combout(\Add1~15_combout ),
	.cout());
defparam \Add1~15 .lut_mask = 16'h0FF0;
defparam \Add1~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[13]~15 (
	.dataa(\D_iw[17]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[13]~15_combout ),
	.cout());
defparam \E_src1[13]~15 .lut_mask = 16'hAACC;
defparam \E_src1[13]~15 .sum_lutc_input = "datac";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\E_src1[13]~15_combout ),
	.asdata(\F_pc_plus_one[11]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[12]~3 (
	.dataa(\D_iw[18]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[12]~3_combout ),
	.cout());
defparam \R_src2_lo[12]~3 .lut_mask = 16'hACFF;
defparam \R_src2_lo[12]~3 .sum_lutc_input = "datac";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\R_src2_lo[12]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cycloneive_lcell_comb \Add1~16 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[12]~q ),
	.cin(gnd),
	.combout(\Add1~16_combout ),
	.cout());
defparam \Add1~16 .lut_mask = 16'h0FF0;
defparam \Add1~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[12]~16 (
	.dataa(\D_iw[16]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[12]~16_combout ),
	.cout());
defparam \E_src1[12]~16 .lut_mask = 16'hAACC;
defparam \E_src1[12]~16 .sum_lutc_input = "datac";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\E_src1[12]~16_combout ),
	.asdata(\F_pc_plus_one[10]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[11]~4 (
	.dataa(\D_iw[17]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[11]~4_combout ),
	.cout());
defparam \R_src2_lo[11]~4 .lut_mask = 16'hACFF;
defparam \R_src2_lo[11]~4 .sum_lutc_input = "datac";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\R_src2_lo[11]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cycloneive_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[11]~q ),
	.cin(gnd),
	.combout(\Add1~17_combout ),
	.cout());
defparam \Add1~17 .lut_mask = 16'h0FF0;
defparam \Add1~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[11]~17 (
	.dataa(\D_iw[15]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[11]~17_combout ),
	.cout());
defparam \E_src1[11]~17 .lut_mask = 16'hAACC;
defparam \E_src1[11]~17 .sum_lutc_input = "datac";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\E_src1[11]~17_combout ),
	.asdata(\F_pc_plus_one[9]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[10]~5 (
	.dataa(\D_iw[16]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[10]~5_combout ),
	.cout());
defparam \R_src2_lo[10]~5 .lut_mask = 16'hACFF;
defparam \R_src2_lo[10]~5 .sum_lutc_input = "datac";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\R_src2_lo[10]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cycloneive_lcell_comb \Add1~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[10]~q ),
	.cin(gnd),
	.combout(\Add1~18_combout ),
	.cout());
defparam \Add1~18 .lut_mask = 16'h0FF0;
defparam \Add1~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[10]~18 (
	.dataa(\D_iw[14]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[10]~18_combout ),
	.cout());
defparam \E_src1[10]~18 .lut_mask = 16'hAACC;
defparam \E_src1[10]~18 .sum_lutc_input = "datac";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\E_src1[10]~18_combout ),
	.asdata(\F_pc_plus_one[8]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[9]~6 (
	.dataa(\D_iw[15]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[9]~6_combout ),
	.cout());
defparam \R_src2_lo[9]~6 .lut_mask = 16'hACFF;
defparam \R_src2_lo[9]~6 .sum_lutc_input = "datac";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\R_src2_lo[9]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cycloneive_lcell_comb \Add1~19 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[9]~q ),
	.cin(gnd),
	.combout(\Add1~19_combout ),
	.cout());
defparam \Add1~19 .lut_mask = 16'h0FF0;
defparam \Add1~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[9]~19 (
	.dataa(\D_iw[13]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[9]~19_combout ),
	.cout());
defparam \E_src1[9]~19 .lut_mask = 16'hAACC;
defparam \E_src1[9]~19 .sum_lutc_input = "datac";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\E_src1[9]~19_combout ),
	.asdata(\F_pc_plus_one[7]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[8]~7 (
	.dataa(\D_iw[14]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[8]~7_combout ),
	.cout());
defparam \R_src2_lo[8]~7 .lut_mask = 16'hACFF;
defparam \R_src2_lo[8]~7 .sum_lutc_input = "datac";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\R_src2_lo[8]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cycloneive_lcell_comb \Add1~20 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[8]~q ),
	.cin(gnd),
	.combout(\Add1~20_combout ),
	.cout());
defparam \Add1~20 .lut_mask = 16'h0FF0;
defparam \Add1~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[8]~20 (
	.dataa(\D_iw[12]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[8]~20_combout ),
	.cout());
defparam \E_src1[8]~20 .lut_mask = 16'hAACC;
defparam \E_src1[8]~20 .sum_lutc_input = "datac";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\E_src1[8]~20_combout ),
	.asdata(\F_pc_plus_one[6]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[7]~8 (
	.dataa(\D_iw[13]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[7]~8_combout ),
	.cout());
defparam \R_src2_lo[7]~8 .lut_mask = 16'hACFF;
defparam \R_src2_lo[7]~8 .sum_lutc_input = "datac";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\R_src2_lo[7]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cycloneive_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[7]~q ),
	.cin(gnd),
	.combout(\Add1~21_combout ),
	.cout());
defparam \Add1~21 .lut_mask = 16'h0FF0;
defparam \Add1~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[7]~21 (
	.dataa(\D_iw[11]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[7]~21_combout ),
	.cout());
defparam \E_src1[7]~21 .lut_mask = 16'hAACC;
defparam \E_src1[7]~21 .sum_lutc_input = "datac";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\E_src1[7]~21_combout ),
	.asdata(\F_pc_plus_one[5]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[6]~9 (
	.dataa(\D_iw[12]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[6]~9_combout ),
	.cout());
defparam \R_src2_lo[6]~9 .lut_mask = 16'hACFF;
defparam \R_src2_lo[6]~9 .sum_lutc_input = "datac";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\R_src2_lo[6]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cycloneive_lcell_comb \Add1~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[6]~q ),
	.cin(gnd),
	.combout(\Add1~22_combout ),
	.cout());
defparam \Add1~22 .lut_mask = 16'h0FF0;
defparam \Add1~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[6]~22 (
	.dataa(\D_iw[10]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[6]~22_combout ),
	.cout());
defparam \E_src1[6]~22 .lut_mask = 16'hAACC;
defparam \E_src1[6]~22 .sum_lutc_input = "datac";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~22_combout ),
	.asdata(\F_pc_plus_one[4]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[5]~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[5]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[5]~10_combout ),
	.cout());
defparam \R_src2_lo[5]~10 .lut_mask = 16'hACFF;
defparam \R_src2_lo[5]~10 .sum_lutc_input = "datac";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\R_src2_lo[5]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cycloneive_lcell_comb \Add1~23 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[5]~q ),
	.cin(gnd),
	.combout(\Add1~23_combout ),
	.cout());
defparam \Add1~23 .lut_mask = 16'h0FF0;
defparam \Add1~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[5]~23 (
	.dataa(\D_iw[9]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[5]~23_combout ),
	.cout());
defparam \E_src1[5]~23 .lut_mask = 16'hAACC;
defparam \E_src1[5]~23 .sum_lutc_input = "datac";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~23_combout ),
	.asdata(\F_pc_plus_one[3]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cycloneive_lcell_comb \Add1~24 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_src2[4]~q ),
	.datad(\E_alu_sub~q ),
	.cin(gnd),
	.combout(\Add1~24_combout ),
	.cout());
defparam \Add1~24 .lut_mask = 16'h0FF0;
defparam \Add1~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[4]~24 (
	.dataa(\D_iw[8]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[4]~24_combout ),
	.cout());
defparam \E_src1[4]~24 .lut_mask = 16'hAACC;
defparam \E_src1[4]~24 .sum_lutc_input = "datac";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\E_src1[4]~24_combout ),
	.asdata(\F_pc_plus_one[2]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cycloneive_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[3]~q ),
	.cin(gnd),
	.combout(\Add1~25_combout ),
	.cout());
defparam \Add1~25 .lut_mask = 16'h0FF0;
defparam \Add1~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[3]~26 (
	.dataa(\D_iw[7]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[3]~26_combout ),
	.cout());
defparam \E_src1[3]~26 .lut_mask = 16'hAACC;
defparam \E_src1[3]~26 .sum_lutc_input = "datac";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\E_src1[3]~26_combout ),
	.asdata(\F_pc_plus_one[1]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cycloneive_lcell_comb \Add1~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[2]~q ),
	.cin(gnd),
	.combout(\Add1~26_combout ),
	.cout());
defparam \Add1~26 .lut_mask = 16'h0FF0;
defparam \Add1~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[2]~25 (
	.dataa(\D_iw[6]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\R_src1~10_combout ),
	.cin(gnd),
	.combout(\E_src1[2]~25_combout ),
	.cout());
defparam \E_src1[2]~25 .lut_mask = 16'hAACC;
defparam \E_src1[2]~25 .sum_lutc_input = "datac";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\E_src1[2]~25_combout ),
	.asdata(\F_pc_plus_one[0]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~11_combout ),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cycloneive_lcell_comb \Add1~27 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[1]~q ),
	.cin(gnd),
	.combout(\Add1~27_combout ),
	.cout());
defparam \Add1~27 .lut_mask = 16'h0FF0;
defparam \Add1~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~28 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[0]~q ),
	.cin(gnd),
	.combout(\Add1~28_combout ),
	.cout());
defparam \Add1~28 .lut_mask = 16'h0FF0;
defparam \Add1~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~30 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add1~30_cout ));
defparam \Add1~30 .lut_mask = 16'h00AA;
defparam \Add1~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~31 (
	.dataa(\Add1~28_combout ),
	.datab(\E_src1[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~30_cout ),
	.combout(\Add1~31_combout ),
	.cout(\Add1~32 ));
defparam \Add1~31 .lut_mask = 16'h967F;
defparam \Add1~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~33 (
	.dataa(\Add1~27_combout ),
	.datab(\E_src1[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~32 ),
	.combout(\Add1~33_combout ),
	.cout(\Add1~34 ));
defparam \Add1~33 .lut_mask = 16'h96EF;
defparam \Add1~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~35 (
	.dataa(\Add1~26_combout ),
	.datab(\E_src1[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~34 ),
	.combout(\Add1~35_combout ),
	.cout(\Add1~36 ));
defparam \Add1~35 .lut_mask = 16'h967F;
defparam \Add1~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~37 (
	.dataa(\Add1~25_combout ),
	.datab(\E_src1[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~36 ),
	.combout(\Add1~37_combout ),
	.cout(\Add1~38 ));
defparam \Add1~37 .lut_mask = 16'h96EF;
defparam \Add1~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~39 (
	.dataa(\Add1~24_combout ),
	.datab(\E_src1[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~38 ),
	.combout(\Add1~39_combout ),
	.cout(\Add1~40 ));
defparam \Add1~39 .lut_mask = 16'h967F;
defparam \Add1~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~41 (
	.dataa(\Add1~23_combout ),
	.datab(\E_src1[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~40 ),
	.combout(\Add1~41_combout ),
	.cout(\Add1~42 ));
defparam \Add1~41 .lut_mask = 16'h96EF;
defparam \Add1~41 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~43 (
	.dataa(\Add1~22_combout ),
	.datab(\E_src1[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~42 ),
	.combout(\Add1~43_combout ),
	.cout(\Add1~44 ));
defparam \Add1~43 .lut_mask = 16'h967F;
defparam \Add1~43 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~45 (
	.dataa(\Add1~21_combout ),
	.datab(\E_src1[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~44 ),
	.combout(\Add1~45_combout ),
	.cout(\Add1~46 ));
defparam \Add1~45 .lut_mask = 16'h96EF;
defparam \Add1~45 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~47 (
	.dataa(\Add1~20_combout ),
	.datab(\E_src1[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~46 ),
	.combout(\Add1~47_combout ),
	.cout(\Add1~48 ));
defparam \Add1~47 .lut_mask = 16'h967F;
defparam \Add1~47 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~49 (
	.dataa(\Add1~19_combout ),
	.datab(\E_src1[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~48 ),
	.combout(\Add1~49_combout ),
	.cout(\Add1~50 ));
defparam \Add1~49 .lut_mask = 16'h96EF;
defparam \Add1~49 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~51 (
	.dataa(\Add1~18_combout ),
	.datab(\E_src1[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~50 ),
	.combout(\Add1~51_combout ),
	.cout(\Add1~52 ));
defparam \Add1~51 .lut_mask = 16'h967F;
defparam \Add1~51 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~53 (
	.dataa(\Add1~17_combout ),
	.datab(\E_src1[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~52 ),
	.combout(\Add1~53_combout ),
	.cout(\Add1~54 ));
defparam \Add1~53 .lut_mask = 16'h96EF;
defparam \Add1~53 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~55 (
	.dataa(\Add1~16_combout ),
	.datab(\E_src1[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~54 ),
	.combout(\Add1~55_combout ),
	.cout(\Add1~56 ));
defparam \Add1~55 .lut_mask = 16'h967F;
defparam \Add1~55 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~57 (
	.dataa(\Add1~15_combout ),
	.datab(\E_src1[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~56 ),
	.combout(\Add1~57_combout ),
	.cout(\Add1~58 ));
defparam \Add1~57 .lut_mask = 16'h96EF;
defparam \Add1~57 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~59 (
	.dataa(\Add1~14_combout ),
	.datab(\E_src1[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~58 ),
	.combout(\Add1~59_combout ),
	.cout(\Add1~60 ));
defparam \Add1~59 .lut_mask = 16'h967F;
defparam \Add1~59 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~61 (
	.dataa(\Add1~13_combout ),
	.datab(\E_src1[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~60 ),
	.combout(\Add1~61_combout ),
	.cout(\Add1~62 ));
defparam \Add1~61 .lut_mask = 16'h96EF;
defparam \Add1~61 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~63 (
	.dataa(\Add1~12_combout ),
	.datab(\E_src1[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~62 ),
	.combout(\Add1~63_combout ),
	.cout(\Add1~64 ));
defparam \Add1~63 .lut_mask = 16'h967F;
defparam \Add1~63 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~65 (
	.dataa(\Add1~11_combout ),
	.datab(\E_src1[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~64 ),
	.combout(\Add1~65_combout ),
	.cout(\Add1~66 ));
defparam \Add1~65 .lut_mask = 16'h96EF;
defparam \Add1~65 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~67 (
	.dataa(\Add1~10_combout ),
	.datab(\E_src1[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~66 ),
	.combout(\Add1~67_combout ),
	.cout(\Add1~68 ));
defparam \Add1~67 .lut_mask = 16'h967F;
defparam \Add1~67 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~69 (
	.dataa(\Add1~9_combout ),
	.datab(\E_src1[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~68 ),
	.combout(\Add1~69_combout ),
	.cout(\Add1~70 ));
defparam \Add1~69 .lut_mask = 16'h96EF;
defparam \Add1~69 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~71 (
	.dataa(\Add1~8_combout ),
	.datab(\E_src1[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~70 ),
	.combout(\Add1~71_combout ),
	.cout(\Add1~72 ));
defparam \Add1~71 .lut_mask = 16'h967F;
defparam \Add1~71 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~73 (
	.dataa(\Add1~7_combout ),
	.datab(\E_src1[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~72 ),
	.combout(\Add1~73_combout ),
	.cout(\Add1~74 ));
defparam \Add1~73 .lut_mask = 16'h96EF;
defparam \Add1~73 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~75 (
	.dataa(\Add1~6_combout ),
	.datab(\E_src1[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~74 ),
	.combout(\Add1~75_combout ),
	.cout(\Add1~76 ));
defparam \Add1~75 .lut_mask = 16'h967F;
defparam \Add1~75 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~77 (
	.dataa(\Add1~5_combout ),
	.datab(\E_src1[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~76 ),
	.combout(\Add1~77_combout ),
	.cout(\Add1~78 ));
defparam \Add1~77 .lut_mask = 16'h96EF;
defparam \Add1~77 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~79 (
	.dataa(\Add1~4_combout ),
	.datab(\E_src1[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~78 ),
	.combout(\Add1~79_combout ),
	.cout(\Add1~80 ));
defparam \Add1~79 .lut_mask = 16'h967F;
defparam \Add1~79 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~81 (
	.dataa(\Add1~3_combout ),
	.datab(\E_src1[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~80 ),
	.combout(\Add1~81_combout ),
	.cout(\Add1~82 ));
defparam \Add1~81 .lut_mask = 16'h96EF;
defparam \Add1~81 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~83 (
	.dataa(\Add1~2_combout ),
	.datab(\E_src1[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~82 ),
	.combout(\Add1~83_combout ),
	.cout(\Add1~84 ));
defparam \Add1~83 .lut_mask = 16'h967F;
defparam \Add1~83 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~85 (
	.dataa(\Add1~1_combout ),
	.datab(\E_src1[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~84 ),
	.combout(\Add1~85_combout ),
	.cout(\Add1~86 ));
defparam \Add1~85 .lut_mask = 16'h96EF;
defparam \Add1~85 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~87 (
	.dataa(\Add1~0_combout ),
	.datab(\E_src1[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~86 ),
	.combout(\Add1~87_combout ),
	.cout(\Add1~88 ));
defparam \Add1~87 .lut_mask = 16'h967F;
defparam \Add1~87 .sum_lutc_input = "cin";

cycloneive_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.cout());
defparam \D_logic_op_raw[1]~0 .lut_mask = 16'hEFFF;
defparam \D_logic_op_raw[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~10 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(\D_ctrl_alu_force_xor~14_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~10_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~10 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~11 (
	.dataa(\Equal0~5_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~11_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~11 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~13 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~13_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~13 .lut_mask = 16'hFFD8;
defparam \D_ctrl_alu_force_xor~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~12 (
	.dataa(\D_ctrl_alu_force_xor~10_combout ),
	.datab(\D_ctrl_alu_force_xor~11_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_force_xor~13_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~12_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~12 .lut_mask = 16'hFFFE;
defparam \D_ctrl_alu_force_xor~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_logic_op[1]~0 (
	.dataa(\D_logic_op_raw[1]~0_combout ),
	.datab(\D_ctrl_alu_force_xor~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.cout());
defparam \D_logic_op[1]~0 .lut_mask = 16'hEEEE;
defparam \D_logic_op[1]~0 .sum_lutc_input = "datac";

dffeas \R_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op[0]~1 (
	.dataa(\D_ctrl_alu_force_xor~12_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\Equal0~7_combout ),
	.cin(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.cout());
defparam \D_logic_op[0]~1 .lut_mask = 16'hFAFC;
defparam \D_logic_op[0]~1 .sum_lutc_input = "datac";

dffeas \R_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[28]~0 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[28]~q ),
	.datac(\E_src1[28]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[28]~0_combout ),
	.cout());
defparam \E_logic_result[28]~0 .lut_mask = 16'h6996;
defparam \E_logic_result[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~8 (
	.dataa(\D_iw[13]~q ),
	.datab(gnd),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'hAFFF;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_ctrl_logic(
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\Equal0~8_combout ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~combout ),
	.cout());
defparam D_ctrl_logic.lut_mask = 16'hFEFF;
defparam D_ctrl_logic.sum_lutc_input = "datac";

dffeas R_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cycloneive_lcell_comb \W_alu_result[28]~0 (
	.dataa(\Add1~87_combout ),
	.datab(\E_logic_result[28]~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[28]~0_combout ),
	.cout());
defparam \W_alu_result[28]~0 .lut_mask = 16'hAACC;
defparam \W_alu_result[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_shift_rot_right~0_combout ),
	.datad(\D_iw[13]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~1 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[27]~1 (
	.dataa(\E_shift_rot_result[28]~q ),
	.datab(\E_shift_rot_result[26]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[27]~1_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[27]~1 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[27]~1 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[27]~1_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[26]~2 (
	.dataa(\E_shift_rot_result[27]~q ),
	.datab(\E_shift_rot_result[25]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[26]~2_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[26]~2 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[26]~2 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[26]~2_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[25]~3 (
	.dataa(\E_shift_rot_result[26]~q ),
	.datab(\E_shift_rot_result[24]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[25]~3_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[25]~3 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[25]~3 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[25]~3_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[24]~4 (
	.dataa(\E_shift_rot_result[25]~q ),
	.datab(\E_shift_rot_result[23]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[24]~4_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[24]~4 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[24]~4 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[24]~4_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[23]~5 (
	.dataa(\E_shift_rot_result[24]~q ),
	.datab(\E_shift_rot_result[22]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[23]~5_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[23]~5 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[23]~5 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[23]~5_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[22]~6 (
	.dataa(\E_shift_rot_result[23]~q ),
	.datab(\E_shift_rot_result[21]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[22]~6_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[22]~6 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[22]~6 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[22]~6_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[21]~7 (
	.dataa(\E_shift_rot_result[22]~q ),
	.datab(\E_shift_rot_result[20]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[21]~7_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[21]~7 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[21]~7 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[21]~7_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[20]~8 (
	.dataa(\E_shift_rot_result[21]~q ),
	.datab(\E_shift_rot_result[19]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[20]~8_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[20]~8 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[20]~8 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[20]~8_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[19]~9 (
	.dataa(\E_shift_rot_result[20]~q ),
	.datab(\E_shift_rot_result[18]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[19]~9_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[19]~9 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[19]~9 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[19]~9_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[18]~10 (
	.dataa(\E_shift_rot_result[19]~q ),
	.datab(\E_shift_rot_result[17]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[18]~10_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[18]~10 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[18]~10 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[18]~10_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[17]~11 (
	.dataa(\E_shift_rot_result[18]~q ),
	.datab(\E_shift_rot_result[16]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[17]~11_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[17]~11 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[17]~11 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[17]~11_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[16]~12 (
	.dataa(\E_shift_rot_result[17]~q ),
	.datab(\E_shift_rot_result[15]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[16]~12_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[16]~12 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[16]~12 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[16]~12_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[15]~13 (
	.dataa(\E_shift_rot_result[16]~q ),
	.datab(\E_shift_rot_result[14]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[15]~13_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[15]~13 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[15]~13 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[15]~13_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[14]~14 (
	.dataa(\E_shift_rot_result[15]~q ),
	.datab(\E_shift_rot_result[13]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[14]~14_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[14]~14 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[14]~14 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[14]~14_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[13]~15 (
	.dataa(\E_shift_rot_result[14]~q ),
	.datab(\E_shift_rot_result[12]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[13]~15_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[13]~15 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[13]~15 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[13]~15_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[12]~20 (
	.dataa(\E_shift_rot_result[13]~q ),
	.datab(\E_shift_rot_result[11]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[12]~20_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[12]~20 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[12]~20 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[12]~20_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[11]~24 (
	.dataa(\E_shift_rot_result[12]~q ),
	.datab(\E_shift_rot_result[10]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[11]~24_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[11]~24 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[11]~24 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[11]~24_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[10]~21 (
	.dataa(\E_shift_rot_result[11]~q ),
	.datab(\E_shift_rot_result[9]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[10]~21_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[10]~21 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[10]~21 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[10]~21_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[9]~22 (
	.dataa(\E_shift_rot_result[10]~q ),
	.datab(\E_shift_rot_result[8]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[9]~22_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[9]~22 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[9]~22 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[9]~22_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[8]~23 (
	.dataa(\E_shift_rot_result[9]~q ),
	.datab(\E_shift_rot_result[7]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[8]~23_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[8]~23 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[8]~23 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[8]~23_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[7]~17 (
	.dataa(\E_shift_rot_result[8]~q ),
	.datab(\E_shift_rot_result[6]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[7]~17_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[7]~17 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[7]~17 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[7]~17_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[6]~16 (
	.dataa(\E_shift_rot_result[7]~q ),
	.datab(\E_shift_rot_result[5]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[6]~16_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[6]~16 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[6]~16 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[6]~16_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[5]~18 (
	.dataa(\E_shift_rot_result[6]~q ),
	.datab(\E_shift_rot_result[4]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[5]~18_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[5]~18 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[5]~18 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[5]~18_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[4]~19 (
	.dataa(\E_shift_rot_result[5]~q ),
	.datab(\E_shift_rot_result[3]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[4]~19_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[4]~19 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[4]~19 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[4]~19_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[3]~26 (
	.dataa(\E_shift_rot_result[4]~q ),
	.datab(\E_shift_rot_result[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[3]~26_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[3]~26 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[3]~26 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[3]~26_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[2]~25 (
	.dataa(\E_shift_rot_result[3]~q ),
	.datab(\E_shift_rot_result[1]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[2]~25_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[2]~25 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[2]~25 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[2]~25_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[1]~28 (
	.dataa(\E_shift_rot_result[2]~q ),
	.datab(\E_shift_rot_result[0]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[1]~28_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[1]~28 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[1]~28 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[1]~28_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[0]~30 (
	.dataa(\E_shift_rot_result[1]~q ),
	.datab(\E_shift_rot_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[0]~30_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[0]~30 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[0]~30 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[0]~30_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cycloneive_lcell_comb \R_ctrl_rot_right_nxt~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~7_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\R_ctrl_rot_right_nxt~0_combout ),
	.cout());
defparam \R_ctrl_rot_right_nxt~0 .lut_mask = 16'hFEFF;
defparam \R_ctrl_rot_right_nxt~0 .sum_lutc_input = "datac";

dffeas R_ctrl_rot_right(
	.clk(clk_clk),
	.d(\R_ctrl_rot_right_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cycloneive_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~4_combout ),
	.datad(\Equal62~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.cout());
defparam \D_ctrl_shift_logical~1 .lut_mask = 16'hFFB8;
defparam \D_ctrl_shift_logical~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[15]~q ),
	.datac(\D_ctrl_shift_logical~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~2_combout ),
	.cout());
defparam \D_ctrl_shift_logical~2 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_logical~2 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(\E_shift_rot_result[0]~q ),
	.datab(\E_shift_rot_result[31]~q ),
	.datac(\R_ctrl_rot_right~q ),
	.datad(\R_ctrl_shift_logical~q ),
	.cin(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.cout());
defparam \E_shift_rot_fill_bit~0 .lut_mask = 16'hACFF;
defparam \E_shift_rot_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_result_nxt[31]~31 (
	.dataa(\E_shift_rot_fill_bit~0_combout ),
	.datab(\E_shift_rot_result[30]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[31]~31_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[31]~31 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[31]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[31]~14 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[31]~14_combout ),
	.cout());
defparam \R_src1[31]~14 .lut_mask = 16'hF7FF;
defparam \R_src1[31]~14 .sum_lutc_input = "datac";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\R_src1[31]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[31]~31_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[30]~29 (
	.dataa(\E_shift_rot_result[31]~q ),
	.datab(\E_shift_rot_result[29]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[30]~29_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[30]~29 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[30]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[30]~15 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[30]~15_combout ),
	.cout());
defparam \R_src1[30]~15 .lut_mask = 16'hF7FF;
defparam \R_src1[30]~15 .sum_lutc_input = "datac";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\R_src1[30]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[30]~29_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[29]~27 (
	.dataa(\E_shift_rot_result[30]~q ),
	.datab(\E_shift_rot_result[28]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[29]~27_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[29]~27 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[29]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[29]~16 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\final_project_soc_nios2_qsys_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(\R_src1~11_combout ),
	.cin(gnd),
	.combout(\R_src1[29]~16_combout ),
	.cout());
defparam \R_src1[29]~16 .lut_mask = 16'hF7FF;
defparam \R_src1[29]~16 .sum_lutc_input = "datac";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\R_src1[29]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[29]~27_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[28]~0 (
	.dataa(\E_shift_rot_result[29]~q ),
	.datab(\E_shift_rot_result[27]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[28]~0_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[28]~0 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[28]~0 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[28]~0_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cycloneive_lcell_comb D_op_rdctl(
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_rdctl~combout ),
	.cout());
defparam D_op_rdctl.lut_mask = 16'hEFFF;
defparam D_op_rdctl.sum_lutc_input = "datac";

dffeas R_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cycloneive_lcell_comb \D_ctrl_br_cmp~2 (
	.dataa(\Equal0~6_combout ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~3_combout ),
	.datad(\D_ctrl_jmp_direct~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~2_combout ),
	.cout());
defparam \D_ctrl_br_cmp~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_br_cmp~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~5 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~5_combout ),
	.cout());
defparam \D_ctrl_br_cmp~5 .lut_mask = 16'hF7B3;
defparam \D_ctrl_br_cmp~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~3 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\D_ctrl_br_cmp~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~3_combout ),
	.cout());
defparam \D_ctrl_br_cmp~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_br_cmp~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~4 (
	.dataa(\D_ctrl_br_cmp~2_combout ),
	.datab(\D_ctrl_br_cmp~3_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~4_combout ),
	.cout());
defparam \D_ctrl_br_cmp~4 .lut_mask = 16'hFFFE;
defparam \D_ctrl_br_cmp~4 .sum_lutc_input = "datac";

dffeas R_ctrl_br_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_br_cmp~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cycloneive_lcell_comb \E_alu_result~0 (
	.dataa(\R_ctrl_rd_ctl_reg~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_alu_result~0_combout ),
	.cout());
defparam \E_alu_result~0 .lut_mask = 16'hEEEE;
defparam \E_alu_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[27]~1 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[27]~q ),
	.datac(\E_src1[27]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[27]~1_combout ),
	.cout());
defparam \E_logic_result[27]~1 .lut_mask = 16'h6996;
defparam \E_logic_result[27]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[27]~1 (
	.dataa(\Add1~85_combout ),
	.datab(\E_logic_result[27]~1_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[27]~1_combout ),
	.cout());
defparam \W_alu_result[27]~1 .lut_mask = 16'hAACC;
defparam \W_alu_result[27]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[26]~2 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[26]~q ),
	.datac(\E_src1[26]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[26]~2_combout ),
	.cout());
defparam \E_logic_result[26]~2 .lut_mask = 16'h6996;
defparam \E_logic_result[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[26]~2 (
	.dataa(\Add1~83_combout ),
	.datab(\E_logic_result[26]~2_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[26]~2_combout ),
	.cout());
defparam \W_alu_result[26]~2 .lut_mask = 16'hAACC;
defparam \W_alu_result[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[25]~3 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[25]~q ),
	.datac(\E_src1[25]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[25]~3_combout ),
	.cout());
defparam \E_logic_result[25]~3 .lut_mask = 16'h6996;
defparam \E_logic_result[25]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[25]~3 (
	.dataa(\Add1~81_combout ),
	.datab(\E_logic_result[25]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[25]~3_combout ),
	.cout());
defparam \W_alu_result[25]~3 .lut_mask = 16'hAACC;
defparam \W_alu_result[25]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[24]~4 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[24]~q ),
	.datac(\E_src1[24]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[24]~4_combout ),
	.cout());
defparam \E_logic_result[24]~4 .lut_mask = 16'h6996;
defparam \E_logic_result[24]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[24]~4 (
	.dataa(\Add1~79_combout ),
	.datab(\E_logic_result[24]~4_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[24]~4_combout ),
	.cout());
defparam \W_alu_result[24]~4 .lut_mask = 16'hAACC;
defparam \W_alu_result[24]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[23]~5 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[23]~q ),
	.datac(\E_src1[23]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[23]~5_combout ),
	.cout());
defparam \E_logic_result[23]~5 .lut_mask = 16'h6996;
defparam \E_logic_result[23]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[23]~5 (
	.dataa(\Add1~77_combout ),
	.datab(\E_logic_result[23]~5_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[23]~5_combout ),
	.cout());
defparam \W_alu_result[23]~5 .lut_mask = 16'hAACC;
defparam \W_alu_result[23]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[22]~6 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[22]~q ),
	.datac(\E_src1[22]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[22]~6_combout ),
	.cout());
defparam \E_logic_result[22]~6 .lut_mask = 16'h6996;
defparam \E_logic_result[22]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[22]~6 (
	.dataa(\Add1~75_combout ),
	.datab(\E_logic_result[22]~6_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[22]~6_combout ),
	.cout());
defparam \W_alu_result[22]~6 .lut_mask = 16'hAACC;
defparam \W_alu_result[22]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[21]~7 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[21]~q ),
	.datac(\E_src1[21]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[21]~7_combout ),
	.cout());
defparam \E_logic_result[21]~7 .lut_mask = 16'h6996;
defparam \E_logic_result[21]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[21]~7 (
	.dataa(\Add1~73_combout ),
	.datab(\E_logic_result[21]~7_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[21]~7_combout ),
	.cout());
defparam \W_alu_result[21]~7 .lut_mask = 16'hAACC;
defparam \W_alu_result[21]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[20]~8 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[20]~q ),
	.datac(\E_src1[20]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[20]~8_combout ),
	.cout());
defparam \E_logic_result[20]~8 .lut_mask = 16'h6996;
defparam \E_logic_result[20]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[20]~8 (
	.dataa(\Add1~71_combout ),
	.datab(\E_logic_result[20]~8_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[20]~8_combout ),
	.cout());
defparam \W_alu_result[20]~8 .lut_mask = 16'hAACC;
defparam \W_alu_result[20]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[19]~9 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[19]~q ),
	.datac(\E_src1[19]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[19]~9_combout ),
	.cout());
defparam \E_logic_result[19]~9 .lut_mask = 16'h6996;
defparam \E_logic_result[19]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[19]~9 (
	.dataa(\Add1~69_combout ),
	.datab(\E_logic_result[19]~9_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[19]~9_combout ),
	.cout());
defparam \W_alu_result[19]~9 .lut_mask = 16'hAACC;
defparam \W_alu_result[19]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[18]~10 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[18]~q ),
	.datac(\E_src1[18]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[18]~10_combout ),
	.cout());
defparam \E_logic_result[18]~10 .lut_mask = 16'h6996;
defparam \E_logic_result[18]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[18]~10 (
	.dataa(\Add1~67_combout ),
	.datab(\E_logic_result[18]~10_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[18]~10_combout ),
	.cout());
defparam \W_alu_result[18]~10 .lut_mask = 16'hAACC;
defparam \W_alu_result[18]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[17]~11 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[17]~q ),
	.datac(\E_src1[17]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[17]~11_combout ),
	.cout());
defparam \E_logic_result[17]~11 .lut_mask = 16'h6996;
defparam \E_logic_result[17]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[17]~11 (
	.dataa(\Add1~65_combout ),
	.datab(\E_logic_result[17]~11_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[17]~11_combout ),
	.cout());
defparam \W_alu_result[17]~11 .lut_mask = 16'hAACC;
defparam \W_alu_result[17]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[16]~12 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[16]~q ),
	.datac(\E_src1[16]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[16]~12_combout ),
	.cout());
defparam \E_logic_result[16]~12 .lut_mask = 16'h6996;
defparam \E_logic_result[16]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[16]~12 (
	.dataa(\Add1~63_combout ),
	.datab(\E_logic_result[16]~12_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[16]~12_combout ),
	.cout());
defparam \W_alu_result[16]~12 .lut_mask = 16'hAACC;
defparam \W_alu_result[16]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[15]~13 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[15]~q ),
	.datac(\E_src1[15]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[15]~13_combout ),
	.cout());
defparam \E_logic_result[15]~13 .lut_mask = 16'h6996;
defparam \E_logic_result[15]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[15]~13 (
	.dataa(\Add1~61_combout ),
	.datab(\E_logic_result[15]~13_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[15]~13_combout ),
	.cout());
defparam \W_alu_result[15]~13 .lut_mask = 16'hAACC;
defparam \W_alu_result[15]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[14]~14 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[14]~q ),
	.datac(\E_src1[14]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[14]~14_combout ),
	.cout());
defparam \E_logic_result[14]~14 .lut_mask = 16'h6996;
defparam \E_logic_result[14]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[14]~14 (
	.dataa(\Add1~59_combout ),
	.datab(\E_logic_result[14]~14_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[14]~14_combout ),
	.cout());
defparam \W_alu_result[14]~14 .lut_mask = 16'hAACC;
defparam \W_alu_result[14]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[13]~15 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[13]~q ),
	.datac(\E_src1[13]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[13]~15_combout ),
	.cout());
defparam \E_logic_result[13]~15 .lut_mask = 16'h6996;
defparam \E_logic_result[13]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[13]~15 (
	.dataa(\Add1~57_combout ),
	.datab(\E_logic_result[13]~15_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[13]~15_combout ),
	.cout());
defparam \W_alu_result[13]~15 .lut_mask = 16'hAACC;
defparam \W_alu_result[13]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[6]~16 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[6]~q ),
	.datac(\E_src1[6]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[6]~16_combout ),
	.cout());
defparam \E_logic_result[6]~16 .lut_mask = 16'h6996;
defparam \E_logic_result[6]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[6]~22 (
	.dataa(\Add1~43_combout ),
	.datab(\E_logic_result[6]~16_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[6]~22_combout ),
	.cout());
defparam \W_alu_result[6]~22 .lut_mask = 16'hAACC;
defparam \W_alu_result[6]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[7]~17 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[7]~q ),
	.datac(\E_src1[7]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[7]~17_combout ),
	.cout());
defparam \E_logic_result[7]~17 .lut_mask = 16'h6996;
defparam \E_logic_result[7]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[7]~21 (
	.dataa(\Add1~45_combout ),
	.datab(\E_logic_result[7]~17_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[7]~21_combout ),
	.cout());
defparam \W_alu_result[7]~21 .lut_mask = 16'hAACC;
defparam \W_alu_result[7]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[5]~18 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[5]~q ),
	.datac(\E_src1[5]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[5]~18_combout ),
	.cout());
defparam \E_logic_result[5]~18 .lut_mask = 16'h6996;
defparam \E_logic_result[5]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[5]~23 (
	.dataa(\Add1~41_combout ),
	.datab(\E_logic_result[5]~18_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[5]~23_combout ),
	.cout());
defparam \W_alu_result[5]~23 .lut_mask = 16'hAACC;
defparam \W_alu_result[5]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[4]~19 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[4]~q ),
	.datac(\E_src1[4]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[4]~19_combout ),
	.cout());
defparam \E_logic_result[4]~19 .lut_mask = 16'h6996;
defparam \E_logic_result[4]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[4]~24 (
	.dataa(\Add1~39_combout ),
	.datab(\E_logic_result[4]~19_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[4]~24_combout ),
	.cout());
defparam \W_alu_result[4]~24 .lut_mask = 16'hAACC;
defparam \W_alu_result[4]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[12]~20 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[12]~q ),
	.datac(\E_src1[12]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[12]~20_combout ),
	.cout());
defparam \E_logic_result[12]~20 .lut_mask = 16'h6996;
defparam \E_logic_result[12]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[12]~16 (
	.dataa(\Add1~55_combout ),
	.datab(\E_logic_result[12]~20_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[12]~16_combout ),
	.cout());
defparam \W_alu_result[12]~16 .lut_mask = 16'hAACC;
defparam \W_alu_result[12]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[10]~21 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[10]~q ),
	.datac(\E_src1[10]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[10]~21_combout ),
	.cout());
defparam \E_logic_result[10]~21 .lut_mask = 16'h6996;
defparam \E_logic_result[10]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[10]~18 (
	.dataa(\Add1~51_combout ),
	.datab(\E_logic_result[10]~21_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[10]~18_combout ),
	.cout());
defparam \W_alu_result[10]~18 .lut_mask = 16'hAACC;
defparam \W_alu_result[10]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[9]~22 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[9]~q ),
	.datac(\E_src1[9]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[9]~22_combout ),
	.cout());
defparam \E_logic_result[9]~22 .lut_mask = 16'h6996;
defparam \E_logic_result[9]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[9]~19 (
	.dataa(\Add1~49_combout ),
	.datab(\E_logic_result[9]~22_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[9]~19_combout ),
	.cout());
defparam \W_alu_result[9]~19 .lut_mask = 16'hAACC;
defparam \W_alu_result[9]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[8]~23 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[8]~q ),
	.datac(\E_src1[8]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[8]~23_combout ),
	.cout());
defparam \E_logic_result[8]~23 .lut_mask = 16'h6996;
defparam \E_logic_result[8]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[8]~20 (
	.dataa(\Add1~47_combout ),
	.datab(\E_logic_result[8]~23_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[8]~20_combout ),
	.cout());
defparam \W_alu_result[8]~20 .lut_mask = 16'hAACC;
defparam \W_alu_result[8]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[11]~24 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[11]~q ),
	.datac(\E_src1[11]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[11]~24_combout ),
	.cout());
defparam \E_logic_result[11]~24 .lut_mask = 16'h6996;
defparam \E_logic_result[11]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[11]~17 (
	.dataa(\Add1~53_combout ),
	.datab(\E_logic_result[11]~24_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[11]~17_combout ),
	.cout());
defparam \W_alu_result[11]~17 .lut_mask = 16'hAACC;
defparam \W_alu_result[11]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[2]~25 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[2]~q ),
	.datac(\E_src1[2]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[2]~25_combout ),
	.cout());
defparam \E_logic_result[2]~25 .lut_mask = 16'h6996;
defparam \E_logic_result[2]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[2]~25 (
	.dataa(\Add1~35_combout ),
	.datab(\E_logic_result[2]~25_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[2]~25_combout ),
	.cout());
defparam \W_alu_result[2]~25 .lut_mask = 16'hAACC;
defparam \W_alu_result[2]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[3]~26 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[3]~q ),
	.datac(\E_src1[3]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[3]~26_combout ),
	.cout());
defparam \E_logic_result[3]~26 .lut_mask = 16'h6996;
defparam \E_logic_result[3]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[3]~26 (
	.dataa(\Add1~37_combout ),
	.datab(\E_logic_result[3]~26_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[3]~26_combout ),
	.cout());
defparam \W_alu_result[3]~26 .lut_mask = 16'hAACC;
defparam \W_alu_result[3]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem16~1 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.cout());
defparam \D_ctrl_mem16~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[31]~3 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[31]~3_combout ),
	.cout());
defparam \d_writedata[31]~3 .lut_mask = 16'hAACC;
defparam \d_writedata[31]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.cout());
defparam \D_ctrl_mem8~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~1 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.cout());
defparam \D_ctrl_mem8~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[30]~4 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[30]~4_combout ),
	.cout());
defparam \d_writedata[30]~4 .lut_mask = 16'hAACC;
defparam \d_writedata[30]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[29]~5 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[29]~5_combout ),
	.cout());
defparam \d_writedata[29]~5 .lut_mask = 16'hAACC;
defparam \d_writedata[29]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[28]~6 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[28]~6_combout ),
	.cout());
defparam \d_writedata[28]~6 .lut_mask = 16'hAACC;
defparam \d_writedata[28]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[27]~7 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[27]~7_combout ),
	.cout());
defparam \d_writedata[27]~7 .lut_mask = 16'hAACC;
defparam \d_writedata[27]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[26]~2 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[26]~2_combout ),
	.cout());
defparam \d_writedata[26]~2 .lut_mask = 16'hAACC;
defparam \d_writedata[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[25]~1 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[25]~1_combout ),
	.cout());
defparam \d_writedata[25]~1 .lut_mask = 16'hAACC;
defparam \d_writedata[25]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[24]~0 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[24]~0_combout ),
	.cout());
defparam \d_writedata[24]~0 .lut_mask = 16'hAACC;
defparam \d_writedata[24]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_read_nxt~0 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(d_read1),
	.datad(av_ld_getting_data),
	.cin(gnd),
	.combout(\d_read_nxt~0_combout ),
	.cout());
defparam \d_read_nxt~0 .lut_mask = 16'hFEFF;
defparam \d_read_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb E_st_stall(
	.dataa(d_write1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_st~q ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\E_st_stall~combout ),
	.cout());
defparam E_st_stall.lut_mask = 16'hFFFE;
defparam E_st_stall.sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~12_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_uncond_cti_non_br~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~2 (
	.dataa(\D_ctrl_jmp_direct~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~2_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~2 .lut_mask = 16'hEEFF;
defparam \D_ctrl_uncond_cti_non_br~2 .sum_lutc_input = "datac";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(clk_clk),
	.d(\D_ctrl_uncond_cti_non_br~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cycloneive_lcell_comb \Equal0~19 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~19_combout ),
	.cout());
defparam \Equal0~19 .lut_mask = 16'hF7F7;
defparam \Equal0~19 .sum_lutc_input = "datac";

dffeas R_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\Equal0~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

dffeas \R_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.cout());
defparam \D_logic_op_raw[0]~1 .lut_mask = 16'hEFFE;
defparam \D_logic_op_raw[0]~1 .sum_lutc_input = "datac";

dffeas \R_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cycloneive_lcell_comb \Equal127~0 (
	.dataa(\E_logic_result[28]~0_combout ),
	.datab(\E_logic_result[27]~1_combout ),
	.datac(\E_logic_result[26]~2_combout ),
	.datad(\E_logic_result[25]~3_combout ),
	.cin(gnd),
	.combout(\Equal127~0_combout ),
	.cout());
defparam \Equal127~0 .lut_mask = 16'h7FFF;
defparam \Equal127~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~1 (
	.dataa(\E_logic_result[24]~4_combout ),
	.datab(\E_logic_result[23]~5_combout ),
	.datac(\E_logic_result[22]~6_combout ),
	.datad(\E_logic_result[21]~7_combout ),
	.cin(gnd),
	.combout(\Equal127~1_combout ),
	.cout());
defparam \Equal127~1 .lut_mask = 16'h7FFF;
defparam \Equal127~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~2 (
	.dataa(\E_logic_result[20]~8_combout ),
	.datab(\E_logic_result[19]~9_combout ),
	.datac(\E_logic_result[18]~10_combout ),
	.datad(\E_logic_result[17]~11_combout ),
	.cin(gnd),
	.combout(\Equal127~2_combout ),
	.cout());
defparam \Equal127~2 .lut_mask = 16'h7FFF;
defparam \Equal127~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~3 (
	.dataa(\E_logic_result[16]~12_combout ),
	.datab(\E_logic_result[15]~13_combout ),
	.datac(\E_logic_result[14]~14_combout ),
	.datad(\E_logic_result[13]~15_combout ),
	.cin(gnd),
	.combout(\Equal127~3_combout ),
	.cout());
defparam \Equal127~3 .lut_mask = 16'h7FFF;
defparam \Equal127~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~4 (
	.dataa(\Equal127~0_combout ),
	.datab(\Equal127~1_combout ),
	.datac(\Equal127~2_combout ),
	.datad(\Equal127~3_combout ),
	.cin(gnd),
	.combout(\Equal127~4_combout ),
	.cout());
defparam \Equal127~4 .lut_mask = 16'hFFFE;
defparam \Equal127~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~5 (
	.dataa(\E_logic_result[11]~24_combout ),
	.datab(\E_logic_result[12]~20_combout ),
	.datac(\E_logic_result[10]~21_combout ),
	.datad(\E_logic_result[9]~22_combout ),
	.cin(gnd),
	.combout(\Equal127~5_combout ),
	.cout());
defparam \Equal127~5 .lut_mask = 16'h7FFF;
defparam \Equal127~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~6 (
	.dataa(\E_logic_result[8]~23_combout ),
	.datab(\E_logic_result[6]~16_combout ),
	.datac(\E_logic_result[7]~17_combout ),
	.datad(\E_logic_result[5]~18_combout ),
	.cin(gnd),
	.combout(\Equal127~6_combout ),
	.cout());
defparam \Equal127~6 .lut_mask = 16'h7FFF;
defparam \Equal127~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~1 (
	.dataa(\D_iw[21]~q ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\R_ctrl_hi_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~1_combout ),
	.cout());
defparam \R_src2_hi[15]~1 .lut_mask = 16'hEFFE;
defparam \R_src2_hi[15]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~2 (
	.dataa(\R_src2_hi[15]~1_combout ),
	.datab(gnd),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(\R_ctrl_unsigned_lo_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~2_combout ),
	.cout());
defparam \R_src2_hi[15]~2 .lut_mask = 16'hAFFF;
defparam \R_src2_hi[15]~2 .sum_lutc_input = "datac";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\R_src2_hi[15]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[31]~27 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_src1[31]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[31]~27_combout ),
	.cout());
defparam \E_logic_result[31]~27 .lut_mask = 16'h6996;
defparam \E_logic_result[31]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~7 (
	.dataa(\E_logic_result[4]~19_combout ),
	.datab(\E_logic_result[2]~25_combout ),
	.datac(\E_logic_result[3]~26_combout ),
	.datad(\E_logic_result[31]~27_combout ),
	.cin(gnd),
	.combout(\Equal127~7_combout ),
	.cout());
defparam \Equal127~7 .lut_mask = 16'h7FFF;
defparam \Equal127~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[30]~13 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[30]~13_combout ),
	.cout());
defparam \E_src2[30]~13 .lut_mask = 16'hAACC;
defparam \E_src2[30]~13 .sum_lutc_input = "datac";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\E_src2[30]~13_combout ),
	.asdata(\D_iw[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[30]~28 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[30]~q ),
	.datac(\E_src1[30]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[30]~28_combout ),
	.cout());
defparam \E_logic_result[30]~28 .lut_mask = 16'h6996;
defparam \E_logic_result[30]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[29]~14 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[29]~14_combout ),
	.cout());
defparam \E_src2[29]~14 .lut_mask = 16'hAACC;
defparam \E_src2[29]~14 .sum_lutc_input = "datac";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\E_src2[29]~14_combout ),
	.asdata(\D_iw[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~0_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[29]~29 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[29]~q ),
	.datac(\E_src1[29]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[29]~29_combout ),
	.cout());
defparam \E_logic_result[29]~29 .lut_mask = 16'h6996;
defparam \E_logic_result[29]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[1]~30 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[1]~q ),
	.datac(\E_src1[1]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[1]~30_combout ),
	.cout());
defparam \E_logic_result[1]~30 .lut_mask = 16'h6996;
defparam \E_logic_result[1]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[0]~31 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[0]~q ),
	.datac(\E_src1[0]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[0]~31_combout ),
	.cout());
defparam \E_logic_result[0]~31 .lut_mask = 16'h6996;
defparam \E_logic_result[0]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~8 (
	.dataa(\E_logic_result[30]~28_combout ),
	.datab(\E_logic_result[29]~29_combout ),
	.datac(\E_logic_result[1]~30_combout ),
	.datad(\E_logic_result[0]~31_combout ),
	.cin(gnd),
	.combout(\Equal127~8_combout ),
	.cout());
defparam \Equal127~8 .lut_mask = 16'h7FFF;
defparam \Equal127~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~9 (
	.dataa(\Equal127~5_combout ),
	.datab(\Equal127~6_combout ),
	.datac(\Equal127~7_combout ),
	.datad(\Equal127~8_combout ),
	.cin(gnd),
	.combout(\Equal127~9_combout ),
	.cout());
defparam \Equal127~9 .lut_mask = 16'hFFFE;
defparam \Equal127~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_cmp_result~0 (
	.dataa(\R_compare_op[1]~q ),
	.datab(\R_compare_op[0]~q ),
	.datac(\Equal127~4_combout ),
	.datad(\Equal127~9_combout ),
	.cin(gnd),
	.combout(\E_cmp_result~0_combout ),
	.cout());
defparam \E_cmp_result~0 .lut_mask = 16'h6996;
defparam \E_cmp_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.cout());
defparam \E_invert_arith_src_msb~0 .lut_mask = 16'hEFFE;
defparam \E_invert_arith_src_msb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(\R_valid~q ),
	.datab(\E_invert_arith_src_msb~0_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_alu_subtract~8_combout ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.cout());
defparam \E_invert_arith_src_msb~1 .lut_mask = 16'hEFFF;
defparam \E_invert_arith_src_msb~1 .sum_lutc_input = "datac";

dffeas E_invert_arith_src_msb(
	.clk(clk_clk),
	.d(\E_invert_arith_src_msb~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cycloneive_lcell_comb \Add1~89 (
	.dataa(\E_alu_sub~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add1~89_combout ),
	.cout());
defparam \Add1~89 .lut_mask = 16'h9696;
defparam \Add1~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_arith_src1[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(\E_src1[31]~q ),
	.cin(gnd),
	.combout(\E_arith_src1[31]~combout ),
	.cout());
defparam \E_arith_src1[31] .lut_mask = 16'h0FF0;
defparam \E_arith_src1[31] .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~90 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[30]~q ),
	.cin(gnd),
	.combout(\Add1~90_combout ),
	.cout());
defparam \Add1~90 .lut_mask = 16'h0FF0;
defparam \Add1~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~91 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[29]~q ),
	.cin(gnd),
	.combout(\Add1~91_combout ),
	.cout());
defparam \Add1~91 .lut_mask = 16'h0FF0;
defparam \Add1~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~98 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~97 ),
	.combout(\Add1~98_combout ),
	.cout());
defparam \Add1~98 .lut_mask = 16'h5A5A;
defparam \Add1~98 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_cmp_result~1 (
	.dataa(\E_cmp_result~0_combout ),
	.datab(\R_compare_op[1]~q ),
	.datac(\Add1~98_combout ),
	.datad(\R_compare_op[0]~q ),
	.cin(gnd),
	.combout(\E_cmp_result~1_combout ),
	.cout());
defparam \E_cmp_result~1 .lut_mask = 16'hEBBE;
defparam \E_cmp_result~1 .sum_lutc_input = "datac";

dffeas W_cmp_result(
	.clk(clk_clk),
	.d(\E_cmp_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cycloneive_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(\R_ctrl_uncond_cti_non_br~q ),
	.datab(\R_ctrl_br_uncond~q ),
	.datac(\W_cmp_result~q ),
	.datad(\R_ctrl_br~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.cout());
defparam \F_pc_sel_nxt~0 .lut_mask = 16'hFFFE;
defparam \F_pc_sel_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[26]~32 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\R_ctrl_break~q ),
	.datad(\F_pc_plus_one[26]~52_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[26]~32_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[26]~32 .lut_mask = 16'hFFDF;
defparam \F_pc_no_crst_nxt[26]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(gnd),
	.datac(\R_ctrl_exception~q ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~0 .lut_mask = 16'hAFFF;
defparam \F_pc_sel_nxt.10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[26]~4 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\F_pc_no_crst_nxt[26]~32_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\Add1~87_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[26]~4_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[26]~4 .lut_mask = 16'h7FFF;
defparam \F_pc_no_crst_nxt[26]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[25]~6 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~85_combout ),
	.datac(\F_pc_plus_one[25]~50_combout ),
	.datad(\F_pc_sel_nxt~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[25]~6_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[25]~6 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[25]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[24]~7 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~83_combout ),
	.datac(\F_pc_plus_one[24]~48_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[24]~7_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[24]~7 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[24]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[23]~8 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~81_combout ),
	.datac(\F_pc_plus_one[23]~46_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[23]~8_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[23]~8 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[23]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[22]~9 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~79_combout ),
	.datac(\F_pc_plus_one[22]~44_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[22]~9_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[22]~9 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[22]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[21]~10 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~77_combout ),
	.datac(\F_pc_plus_one[21]~42_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[21]~10_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[21]~10 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[21]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[20]~11 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~75_combout ),
	.datac(\F_pc_plus_one[20]~40_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[20]~11_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[20]~11 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[20]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[19]~12 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~73_combout ),
	.datac(\F_pc_plus_one[19]~38_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[19]~12_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[19]~12 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[19]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[18]~13 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~71_combout ),
	.datac(\F_pc_plus_one[18]~36_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[18]~13_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[18]~13 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[18]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[17]~14 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~69_combout ),
	.datac(\F_pc_plus_one[17]~34_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[17]~14_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[17]~14 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[17]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[16]~15 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~67_combout ),
	.datac(\F_pc_plus_one[16]~32_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[16]~15_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[16]~15 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[16]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[15]~16 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~65_combout ),
	.datac(\F_pc_plus_one[15]~30_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[15]~16_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[15]~16 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[15]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[14]~17 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~63_combout ),
	.datac(\F_pc_plus_one[14]~28_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[14]~17_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[14]~17 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[14]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[13]~18 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~61_combout ),
	.datac(\F_pc_plus_one[13]~26_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~18_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~18 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[13]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[12]~19 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~59_combout ),
	.datac(\F_pc_plus_one[12]~24_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[12]~19_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[12]~19 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[12]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[11]~20 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~57_combout ),
	.datac(\F_pc_plus_one[11]~22_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[11]~20_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[11]~20 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[11]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[10]~33 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\R_ctrl_exception~q ),
	.datac(\R_ctrl_break~q ),
	.datad(\F_pc_plus_one[10]~20_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~33_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~33 .lut_mask = 16'hFFFD;
defparam \F_pc_no_crst_nxt[10]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[10]~21 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\Add1~55_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_no_crst_nxt[10]~33_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~21_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~21 .lut_mask = 16'hFFFD;
defparam \F_pc_no_crst_nxt[10]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[8]~22 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~51_combout ),
	.datac(\F_pc_plus_one[8]~16_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[8]~22_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[8]~22 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[8]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[7]~23 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~49_combout ),
	.datac(\F_pc_plus_one[7]~14_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[7]~23_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[7]~23 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[7]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[6]~24 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~47_combout ),
	.datac(\F_pc_plus_one[6]~12_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[6]~24_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[6]~24 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[6]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[5]~25 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~45_combout ),
	.datac(\F_pc_plus_one[5]~10_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[5]~25_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[5]~25 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[3]~26 (
	.dataa(\Add1~41_combout ),
	.datab(\F_pc_plus_one[3]~6_combout ),
	.datac(\F_pc_sel_nxt.10~0_combout ),
	.datad(\F_pc_no_crst_nxt[25]~5_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[3]~26_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[3]~26 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[3]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_read_nxt~0 (
	.dataa(\W_valid~q ),
	.datab(gnd),
	.datac(i_read1),
	.datad(av_readdatavalid),
	.cin(gnd),
	.combout(\i_read_nxt~0_combout ),
	.cout());
defparam \i_read_nxt~0 .lut_mask = 16'hFFF5;
defparam \i_read_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[2]~27 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~39_combout ),
	.datac(\F_pc_plus_one[2]~4_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[2]~27_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[2]~27 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[2]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[4]~28 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~43_combout ),
	.datac(\F_pc_plus_one[4]~8_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[4]~28_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[4]~28 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[4]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~29 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~53_combout ),
	.datac(\F_pc_plus_one[9]~18_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~29_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~29 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[9]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[0]~0 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~31_combout ),
	.datad(\Add1~33_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[0]~0_combout ),
	.cout());
defparam \E_mem_byte_en[0]~0 .lut_mask = 16'h6FFF;
defparam \E_mem_byte_en[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[0]~30 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~35_combout ),
	.datac(\F_pc_plus_one[0]~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[0]~30_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[0]~30 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[0]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[1]~31 (
	.dataa(\F_pc_no_crst_nxt[25]~5_combout ),
	.datab(\Add1~37_combout ),
	.datac(\F_pc_plus_one[1]~2_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[1]~31_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[1]~31 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[1]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[8]~0 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[8]~0_combout ),
	.cout());
defparam \E_st_data[8]~0 .lut_mask = 16'hEFFE;
defparam \E_st_data[8]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[9]~1 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[9]~1_combout ),
	.cout());
defparam \E_st_data[9]~1 .lut_mask = 16'hEFFE;
defparam \E_st_data[9]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[10]~2 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[10]~2_combout ),
	.cout());
defparam \E_st_data[10]~2 .lut_mask = 16'hEFFE;
defparam \E_st_data[10]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[11]~3 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[11]~3_combout ),
	.cout());
defparam \E_st_data[11]~3 .lut_mask = 16'hEFFE;
defparam \E_st_data[11]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[12]~4 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[12]~4_combout ),
	.cout());
defparam \E_st_data[12]~4 .lut_mask = 16'hEFFE;
defparam \E_st_data[12]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[13]~5 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[13]~5_combout ),
	.cout());
defparam \E_st_data[13]~5 .lut_mask = 16'hEFFE;
defparam \E_st_data[13]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[14]~6 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[14]~6_combout ),
	.cout());
defparam \E_st_data[14]~6 .lut_mask = 16'hEFFE;
defparam \E_st_data[14]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[15]~7 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[15]~7_combout ),
	.cout());
defparam \E_st_data[15]~7 .lut_mask = 16'hEFFE;
defparam \E_st_data[15]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[22]~8 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(\D_ctrl_mem16~0_combout ),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\d_writedata[22]~8_combout ),
	.cout());
defparam \d_writedata[22]~8 .lut_mask = 16'hEEFF;
defparam \d_writedata[22]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[16]~8 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[16]~8_combout ),
	.cout());
defparam \E_st_data[16]~8 .lut_mask = 16'hAACC;
defparam \E_st_data[16]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[17]~9 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[17]~9_combout ),
	.cout());
defparam \E_st_data[17]~9 .lut_mask = 16'hAACC;
defparam \E_st_data[17]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \hbreak_enabled~0 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~10_combout ),
	.datac(hbreak_enabled1),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.cout());
defparam \hbreak_enabled~0 .lut_mask = 16'hFFF7;
defparam \hbreak_enabled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~33_combout ),
	.datac(\D_ctrl_mem8~1_combout ),
	.datad(\Add1~31_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.cout());
defparam \E_mem_byte_en[2]~1 .lut_mask = 16'hDEFF;
defparam \E_mem_byte_en[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[1]~2 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~31_combout ),
	.datad(\Add1~33_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[1]~2_combout ),
	.cout());
defparam \E_mem_byte_en[1]~2 .lut_mask = 16'hF6FF;
defparam \E_mem_byte_en[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~33_combout ),
	.datac(\Add1~31_combout ),
	.datad(\D_ctrl_mem8~1_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.cout());
defparam \E_mem_byte_en[3]~3 .lut_mask = 16'hFDFE;
defparam \E_mem_byte_en[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[21]~10 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[21]~10_combout ),
	.cout());
defparam \E_st_data[21]~10 .lut_mask = 16'hAACC;
defparam \E_st_data[21]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[18]~11 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[18]~11_combout ),
	.cout());
defparam \E_st_data[18]~11 .lut_mask = 16'hAACC;
defparam \E_st_data[18]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[23]~12 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[23]~12_combout ),
	.cout());
defparam \E_st_data[23]~12 .lut_mask = 16'hAACC;
defparam \E_st_data[23]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[22]~13 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[22]~13_combout ),
	.cout());
defparam \E_st_data[22]~13 .lut_mask = 16'hAACC;
defparam \E_st_data[22]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[20]~14 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[20]~14_combout ),
	.cout());
defparam \E_st_data[20]~14 .lut_mask = 16'hAACC;
defparam \E_st_data[20]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[19]~15 (
	.dataa(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(\final_project_soc_nios2_qsys_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\d_writedata[22]~8_combout ),
	.cin(gnd),
	.combout(\E_st_data[19]~15_combout ),
	.cout());
defparam \E_st_data[19]~15 .lut_mask = 16'hAACC;
defparam \E_st_data[19]~15 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_oci (
	sr_0,
	jtag_break,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	waitrequest,
	mem_used_1,
	WideOr1,
	local_read,
	hbreak_enabled,
	mem,
	address_nxt,
	oci_ienable_1,
	oci_ienable_0,
	oci_single_step_mode,
	r_early_rst,
	readdata_4,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_14,
	readdata_15,
	readdata_21,
	readdata_18,
	readdata_17,
	readdata_31,
	readdata_30,
	readdata_29,
	readdata_28,
	readdata_27,
	readdata_26,
	readdata_25,
	readdata_10,
	readdata_24,
	readdata_9,
	readdata_23,
	readdata_8,
	readdata_22,
	readdata_7,
	readdata_6,
	readdata_20,
	readdata_19,
	debugaccess_nxt,
	writedata_nxt,
	byteenable_nxt,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	jtag_break;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
output 	waitrequest;
input 	mem_used_1;
input 	WideOr1;
input 	local_read;
input 	hbreak_enabled;
input 	mem;
input 	[8:0] address_nxt;
output 	oci_ienable_1;
output 	oci_ienable_0;
output 	oci_single_step_mode;
input 	r_early_rst;
output 	readdata_4;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_14;
output 	readdata_15;
output 	readdata_21;
output 	readdata_18;
output 	readdata_17;
output 	readdata_31;
output 	readdata_30;
output 	readdata_29;
output 	readdata_28;
output 	readdata_27;
output 	readdata_26;
output 	readdata_25;
output 	readdata_10;
output 	readdata_24;
output 	readdata_9;
output 	readdata_23;
output 	readdata_8;
output 	readdata_22;
output 	readdata_7;
output 	readdata_6;
output 	readdata_20;
output 	readdata_19;
input 	debugaccess_nxt;
input 	[31:0] writedata_nxt;
input 	[3:0] byteenable_nxt;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_no_action_break_a~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_ready~q ;
wire \write~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \read~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \debugaccess~q ;
wire \writedata[0]~q ;
wire \address[0]~q ;
wire \address[1]~q ;
wire \address[2]~q ;
wire \address[3]~q ;
wire \address[4]~q ;
wire \address[5]~q ;
wire \address[6]~q ;
wire \address[7]~q ;
wire \byteenable[0]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal0~2_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \writedata[1]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \writedata[3]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \writedata[2]~q ;
wire \writedata[4]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \writedata[13]~q ;
wire \writedata[16]~q ;
wire \byteenable[2]~q ;
wire \writedata[12]~q ;
wire \writedata[5]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \writedata[14]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \writedata[21]~q ;
wire \writedata[18]~q ;
wire \writedata[17]~q ;
wire \writedata[31]~q ;
wire \byteenable[3]~q ;
wire \writedata[30]~q ;
wire \writedata[29]~q ;
wire \writedata[28]~q ;
wire \writedata[27]~q ;
wire \writedata[26]~q ;
wire \writedata[25]~q ;
wire \writedata[10]~q ;
wire \writedata[24]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \writedata[9]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \writedata[23]~q ;
wire \writedata[8]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \writedata[22]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \writedata[7]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \writedata[6]~q ;
wire \writedata[20]~q ;
wire \writedata[19]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \readdata~0_combout ;
wire \address[8]~q ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \readdata~8_combout ;
wire \readdata~9_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~15_combout ;
wire \readdata~16_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;
wire \readdata~20_combout ;
wire \readdata~21_combout ;
wire \readdata~22_combout ;
wire \readdata~23_combout ;
wire \readdata~24_combout ;
wire \readdata~25_combout ;
wire \readdata~26_combout ;
wire \readdata~27_combout ;
wire \readdata~28_combout ;
wire \readdata~29_combout ;
wire \readdata~30_combout ;
wire \readdata~31_combout ;


final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break(
	.break_readreg_0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[1]~q ),
	.jdo_0(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_37(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[37]~q ),
	.jdo_36(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[36]~q ),
	.take_no_action_break_a(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_no_action_break_a~0_combout ),
	.jdo_3(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_17(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_21(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.break_readreg_2(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_31(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_19(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_3(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.break_readreg_16(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_20(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[19]~q ),
	.jdo_23(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_4(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_24(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_17(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.break_readreg_31(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_30(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_29(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_18(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[21]~q ),
	.jdo_22(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_7(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.break_readreg_5(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_24(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_14(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_22(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_6(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[8]~q ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug(
	.jtag_break1(jtag_break),
	.r_sync_rst(r_sync_rst),
	.jdo_35(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.monitor_ready1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_34(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_21(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_25(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_19(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_error1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_error~q ),
	.monitor_go1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_go~q ),
	.jdo_23(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.resetlatch1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_24(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper(
	.sr_0(sr_0),
	.MonDReg_0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[0]~q ),
	.MonDReg_2(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[2]~q ),
	.MonDReg_3(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[3]~q ),
	.MonDReg_4(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_29(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_28(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_11(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_18(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_10(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_8(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[8]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.break_readreg_0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[0]~q ),
	.hbreak_enabled(hbreak_enabled),
	.break_readreg_1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_37(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[37]~q ),
	.jdo_36(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[36]~q ),
	.take_no_action_break_a(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_no_action_break_a~0_combout ),
	.jdo_3(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_35(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.monitor_ready(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_17(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_34(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_21(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.break_readreg_2(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_25(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_33(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_19(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_error(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_error~q ),
	.break_readreg_3(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.break_readreg_16(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_20(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[19]~q ),
	.jdo_23(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_4(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_25(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_27(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_26(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_24(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_17(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[17]~q ),
	.jdo_16(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.resetlatch(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|resetlatch~q ),
	.break_readreg_31(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_30(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[30]~q ),
	.MonDReg_30(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_29(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_13(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_15(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_21(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[21]~q ),
	.MonDReg_9(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_23(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_22(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_7(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[6]~q ),
	.break_readreg_18(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[21]~q ),
	.jdo_22(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_7(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.break_readreg_5(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_24(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_14(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_22(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_6(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break|break_readreg[8]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem(
	.MonDReg_0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[0]~q ),
	.q_a_0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.MonDReg_2(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[2]~q ),
	.q_a_1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.MonDReg_3(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[3]~q ),
	.q_a_11(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_5(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_14(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_21(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_31(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_30(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_29(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_28(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_27(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_26(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_10(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_24(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_9(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_23(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_8(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_22(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_7(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_20(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.MonDReg_4(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_29(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_28(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_11(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_12(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_18(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_10(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_8(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[8]~q ),
	.waitrequest1(waitrequest),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.MonDReg_1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_35(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_17(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_34(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_21(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.r_early_rst(r_early_rst),
	.jdo_4(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.debugaccess(\debugaccess~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_25(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_33(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_19(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.writedata_3(\writedata[3]~q ),
	.jdo_5(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.MonDReg_16(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_20(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[19]~q ),
	.jdo_23(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.writedata_2(\writedata[2]~q ),
	.writedata_4(\writedata[4]~q ),
	.jdo_6(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.MonDReg_25(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_27(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_26(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_24(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_17(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[17]~q ),
	.jdo_16(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_31(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_30(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[30]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.MonDReg_13(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[13]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_16(\writedata[16]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_12(\writedata[12]~q ),
	.writedata_5(\writedata[5]~q ),
	.MonDReg_14(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[14]~q ),
	.writedata_14(\writedata[14]~q ),
	.MonDReg_15(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.MonDReg_21(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[21]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_17(\writedata[17]~q ),
	.writedata_31(\writedata[31]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_10(\writedata[10]~q ),
	.writedata_24(\writedata[24]~q ),
	.MonDReg_9(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[9]~q ),
	.writedata_9(\writedata[9]~q ),
	.MonDReg_23(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[23]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_8(\writedata[8]~q ),
	.MonDReg_22(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[22]~q ),
	.writedata_22(\writedata[22]~q ),
	.MonDReg_7(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[7]~q ),
	.writedata_7(\writedata[7]~q ),
	.MonDReg_6(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|MonDReg[6]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_19(\writedata[19]~q ),
	.jdo_22(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_7(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_14(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper|the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.oci_ienable_1(oci_ienable_1),
	.oci_ienable_0(oci_ienable_0),
	.oci_single_step_mode1(oci_single_step_mode),
	.debugaccess(\debugaccess~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.Equal0(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.take_action_ocireg(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.writedata_1(\writedata[1]~q ),
	.Equal1(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.writedata_3(\writedata[3]~q ),
	.oci_ienable_16(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(waitrequest),
	.datab(WideOr1),
	.datac(mem),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFAFC;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(waitrequest),
	.datab(\read~q ),
	.datac(local_read),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hB8FF;
defparam \read~0 .sum_lutc_input = "datac";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\readdata~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\readdata~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\readdata~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\readdata~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\readdata~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\readdata~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\readdata~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\readdata~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\readdata~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\readdata~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\readdata~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\readdata~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_error~q ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datad(oci_ienable_0),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hB8FF;
defparam \readdata~0 .sum_lutc_input = "datac";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cycloneive_lcell_comb \readdata~1 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datad(oci_ienable_1),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hB8FF;
defparam \readdata~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug|monitor_go~q ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datad(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hFAFC;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~3 (
	.dataa(oci_single_step_mode),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datad(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hFAFC;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hFAFC;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hFAFC;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hFAFC;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hFAFC;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hFAFC;
defparam \readdata~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hFAFC;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~10 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hFAFC;
defparam \readdata~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hFAFC;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hFAFC;
defparam \readdata~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hFAFC;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hFAFC;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hFAFC;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hFAFC;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hFAFC;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hFAFC;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hFAFC;
defparam \readdata~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~20 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hFAFC;
defparam \readdata~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~21 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hFAFC;
defparam \readdata~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~22 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~22_combout ),
	.cout());
defparam \readdata~22 .lut_mask = 16'hFAFC;
defparam \readdata~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~23 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~23_combout ),
	.cout());
defparam \readdata~23 .lut_mask = 16'hFAFC;
defparam \readdata~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~24 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~24_combout ),
	.cout());
defparam \readdata~24 .lut_mask = 16'hFAFC;
defparam \readdata~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~25 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~25_combout ),
	.cout());
defparam \readdata~25 .lut_mask = 16'hFAFC;
defparam \readdata~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~26 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~26_combout ),
	.cout());
defparam \readdata~26 .lut_mask = 16'hFAFC;
defparam \readdata~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~27 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hFAFC;
defparam \readdata~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~28 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hFAFC;
defparam \readdata~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~29 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~29_combout ),
	.cout());
defparam \readdata~29 .lut_mask = 16'hFAFC;
defparam \readdata~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~30 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hFAFC;
defparam \readdata~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~31 (
	.dataa(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~31_combout ),
	.cout());
defparam \readdata~31 .lut_mask = 16'hFAFC;
defparam \readdata~31 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_debug_slave_wrapper (
	sr_0,
	MonDReg_0,
	MonDReg_2,
	MonDReg_3,
	MonDReg_4,
	MonDReg_29,
	MonDReg_28,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_18,
	MonDReg_10,
	MonDReg_8,
	ir_out_0,
	ir_out_1,
	break_readreg_0,
	hbreak_enabled,
	break_readreg_1,
	MonDReg_1,
	jdo_0,
	jdo_37,
	jdo_36,
	take_no_action_break_a,
	jdo_3,
	jdo_35,
	take_action_ocimem_b,
	take_action_ocimem_a,
	monitor_ready,
	jdo_17,
	jdo_34,
	jdo_21,
	jdo_20,
	take_action_ocimem_a1,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_19,
	jdo_18,
	monitor_error,
	break_readreg_3,
	jdo_2,
	jdo_5,
	break_readreg_16,
	MonDReg_16,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	jdo_23,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	MonDReg_26,
	break_readreg_24,
	MonDReg_24,
	break_readreg_17,
	MonDReg_17,
	jdo_16,
	resetlatch,
	break_readreg_31,
	MonDReg_31,
	break_readreg_30,
	MonDReg_30,
	break_readreg_29,
	break_readreg_28,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_21,
	MonDReg_9,
	MonDReg_23,
	MonDReg_22,
	MonDReg_7,
	MonDReg_6,
	break_readreg_18,
	break_readreg_21,
	jdo_22,
	jdo_7,
	break_readreg_5,
	jdo_24,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_22,
	break_readreg_6,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
input 	MonDReg_2;
input 	MonDReg_3;
input 	MonDReg_4;
input 	MonDReg_29;
input 	MonDReg_28;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_18;
input 	MonDReg_10;
input 	MonDReg_8;
output 	ir_out_0;
output 	ir_out_1;
input 	break_readreg_0;
input 	hbreak_enabled;
input 	break_readreg_1;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_37;
output 	jdo_36;
output 	take_no_action_break_a;
output 	jdo_3;
output 	jdo_35;
output 	take_action_ocimem_b;
output 	take_action_ocimem_a;
input 	monitor_ready;
output 	jdo_17;
output 	jdo_34;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a1;
input 	break_readreg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
output 	jdo_19;
output 	jdo_18;
input 	monitor_error;
input 	break_readreg_3;
output 	jdo_2;
output 	jdo_5;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	jdo_23;
input 	break_readreg_4;
output 	jdo_6;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_17;
input 	MonDReg_17;
output 	jdo_16;
input 	resetlatch;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_21;
input 	MonDReg_9;
input 	MonDReg_23;
input 	MonDReg_22;
input 	MonDReg_7;
input 	MonDReg_6;
input 	break_readreg_18;
input 	break_readreg_21;
output 	jdo_22;
output 	jdo_7;
input 	break_readreg_5;
output 	jdo_24;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	break_readreg_22;
input 	break_readreg_6;
input 	break_readreg_15;
input 	break_readreg_23;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[35]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[31]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[7]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[15]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[1]~q ;
wire \final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[2]~q ;
wire \final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[3]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[4]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[37]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[36]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[17]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[34]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[21]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[20]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[5]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[26]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[28]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[27]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[25]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[18]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[33]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[32]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[30]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[29]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[19]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[22]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[6]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[23]~q ;
wire \final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[16]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[24]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[8]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[14]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[13]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[12]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[11]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[10]~q ;
wire \the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[9]~q ;


final_project_soc_sld_virtual_jtag_basic_1 final_project_soc_nios2_qsys_0_cpu_debug_slave_phy(
	.virtual_state_cdr1(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.virtual_state_udr(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk the_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk(
	.sr_0(sr_0),
	.sr_35(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[31]~q ),
	.sr_7(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[15]~q ),
	.sr_1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[2]~q ),
	.virtual_state_uir(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[3]~q ),
	.jdo_0(jdo_0),
	.jdo_37(jdo_37),
	.jdo_36(jdo_36),
	.take_no_action_break_a(take_no_action_break_a),
	.jdo_3(jdo_3),
	.jdo_35(jdo_35),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_17(jdo_17),
	.jdo_34(jdo_34),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.sr_4(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[4]~q ),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_37(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[37]~q ),
	.sr_36(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[36]~q ),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_25(jdo_25),
	.sr_17(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[17]~q ),
	.jdo_33(jdo_33),
	.jdo_32(jdo_32),
	.jdo_31(jdo_31),
	.jdo_30(jdo_30),
	.jdo_29(jdo_29),
	.sr_34(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[34]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.sr_21(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[20]~q ),
	.sr_5(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[5]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.sr_26(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[25]~q ),
	.sr_18(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[18]~q ),
	.sr_33(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[29]~q ),
	.sr_19(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[22]~q ),
	.jdo_23(jdo_23),
	.sr_6(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[6]~q ),
	.jdo_6(jdo_6),
	.jdo_16(jdo_16),
	.sr_23(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[23]~q ),
	.jdo_22(jdo_22),
	.jdo_7(jdo_7),
	.virtual_state_udr(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_24(jdo_24),
	.sr_16(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[16]~q ),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_8(jdo_8),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_11(jdo_11),
	.jdo_10(jdo_10),
	.jdo_9(jdo_9),
	.sr_24(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[24]~q ),
	.sr_8(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[8]~q ),
	.sr_14(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[9]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

final_project_soc_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck(
	.sr_0(sr_0),
	.MonDReg_0(MonDReg_0),
	.MonDReg_2(MonDReg_2),
	.sr_35(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[35]~q ),
	.MonDReg_3(MonDReg_3),
	.sr_31(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[31]~q ),
	.MonDReg_4(MonDReg_4),
	.MonDReg_29(MonDReg_29),
	.MonDReg_28(MonDReg_28),
	.MonDReg_11(MonDReg_11),
	.MonDReg_12(MonDReg_12),
	.MonDReg_5(MonDReg_5),
	.MonDReg_18(MonDReg_18),
	.MonDReg_10(MonDReg_10),
	.MonDReg_8(MonDReg_8),
	.sr_7(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[15]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.sr_1(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[1]~q ),
	.virtual_state_cdr(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.sr_2(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.virtual_state_uir(\final_project_soc_nios2_qsys_0_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.hbreak_enabled(hbreak_enabled),
	.sr_3(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.monitor_ready(monitor_ready),
	.sr_4(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.sr_37(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[37]~q ),
	.sr_36(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[36]~q ),
	.sr_17(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[17]~q ),
	.sr_34(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[34]~q ),
	.sr_21(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[20]~q ),
	.monitor_error(monitor_error),
	.sr_5(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_26(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[27]~q ),
	.sr_25(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[25]~q ),
	.sr_18(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.sr_33(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[29]~q ),
	.sr_19(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_6(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.resetlatch(resetlatch),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.break_readreg_30(break_readreg_30),
	.MonDReg_30(MonDReg_30),
	.break_readreg_29(break_readreg_29),
	.break_readreg_28(break_readreg_28),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.MonDReg_15(MonDReg_15),
	.MonDReg_21(MonDReg_21),
	.MonDReg_9(MonDReg_9),
	.MonDReg_23(MonDReg_23),
	.MonDReg_22(MonDReg_22),
	.MonDReg_7(MonDReg_7),
	.MonDReg_6(MonDReg_6),
	.break_readreg_18(break_readreg_18),
	.sr_23(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.break_readreg_5(break_readreg_5),
	.sr_16(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[16]~q ),
	.sr_24(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.break_readreg_6(break_readreg_6),
	.sr_8(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[8]~q ),
	.break_readreg_15(break_readreg_15),
	.sr_14(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_23(break_readreg_23),
	.break_readreg_7(break_readreg_7),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_10(break_readreg_10),
	.break_readreg_9(break_readreg_9),
	.break_readreg_8(break_readreg_8),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_debug_slave_sysclk (
	sr_0,
	sr_35,
	sr_31,
	sr_7,
	sr_15,
	sr_1,
	sr_2,
	virtual_state_uir,
	sr_3,
	jdo_0,
	jdo_37,
	jdo_36,
	take_no_action_break_a,
	jdo_3,
	jdo_35,
	take_action_ocimem_b1,
	take_action_ocimem_a1,
	jdo_17,
	jdo_34,
	jdo_21,
	jdo_20,
	take_action_ocimem_a2,
	sr_4,
	jdo_1,
	jdo_4,
	sr_37,
	sr_36,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	sr_17,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	sr_34,
	jdo_19,
	jdo_18,
	sr_21,
	sr_20,
	sr_5,
	jdo_2,
	jdo_5,
	sr_26,
	sr_28,
	sr_27,
	sr_25,
	sr_18,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_19,
	sr_22,
	jdo_23,
	sr_6,
	jdo_6,
	jdo_16,
	sr_23,
	jdo_22,
	jdo_7,
	virtual_state_udr,
	jdo_24,
	sr_16,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	sr_24,
	sr_8,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_0;
input 	sr_35;
input 	sr_31;
input 	sr_7;
input 	sr_15;
input 	sr_1;
input 	sr_2;
input 	virtual_state_uir;
input 	sr_3;
output 	jdo_0;
output 	jdo_37;
output 	jdo_36;
output 	take_no_action_break_a;
output 	jdo_3;
output 	jdo_35;
output 	take_action_ocimem_b1;
output 	take_action_ocimem_a1;
output 	jdo_17;
output 	jdo_34;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a2;
input 	sr_4;
output 	jdo_1;
output 	jdo_4;
input 	sr_37;
input 	sr_36;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_25;
input 	sr_17;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
input 	sr_34;
output 	jdo_19;
output 	jdo_18;
input 	sr_21;
input 	sr_20;
input 	sr_5;
output 	jdo_2;
output 	jdo_5;
input 	sr_26;
input 	sr_28;
input 	sr_27;
input 	sr_25;
input 	sr_18;
input 	sr_33;
input 	sr_32;
input 	sr_30;
input 	sr_29;
input 	sr_19;
input 	sr_22;
output 	jdo_23;
input 	sr_6;
output 	jdo_6;
output 	jdo_16;
input 	sr_23;
output 	jdo_22;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_24;
input 	sr_16;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	sr_24;
input 	sr_8;
input 	sr_14;
input 	sr_13;
input 	sr_12;
input 	sr_11;
input 	sr_10;
input 	sr_9;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;
wire \ir[1]~q ;
wire \enable_action_strobe~q ;
wire \ir[0]~q ;


final_project_soc_altera_std_synchronizer_18 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

final_project_soc_altera_std_synchronizer_17 the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

cycloneive_lcell_comb \take_no_action_break_a~0 (
	.dataa(\ir[1]~q ),
	.datab(\enable_action_strobe~q ),
	.datac(gnd),
	.datad(\ir[0]~q ),
	.cin(gnd),
	.combout(take_no_action_break_a),
	.cout());
defparam \take_no_action_break_a~0 .lut_mask = 16'hEEFF;
defparam \take_no_action_break_a~0 .sum_lutc_input = "datac";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_b(
	.dataa(\enable_action_strobe~q ),
	.datab(jdo_35),
	.datac(\ir[1]~q ),
	.datad(\ir[0]~q ),
	.cin(gnd),
	.combout(take_action_ocimem_b1),
	.cout());
defparam take_action_ocimem_b.lut_mask = 16'hEFFF;
defparam take_action_ocimem_b.sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocimem_a~0 (
	.dataa(\enable_action_strobe~q ),
	.datab(gnd),
	.datac(\ir[1]~q ),
	.datad(\ir[0]~q ),
	.cin(gnd),
	.combout(take_action_ocimem_a1),
	.cout());
defparam \take_action_ocimem_a~0 .lut_mask = 16'hAFFF;
defparam \take_action_ocimem_a~0 .sum_lutc_input = "datac";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_a(
	.dataa(jdo_35),
	.datab(gnd),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(take_action_ocimem_a2),
	.cout());
defparam take_action_ocimem_a.lut_mask = 16'hFFF5;
defparam take_action_ocimem_a.sum_lutc_input = "datac";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cycloneive_lcell_comb \update_jdo_strobe~0 (
	.dataa(\the_altera_std_synchronizer3|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_udr~q ),
	.cin(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.cout());
defparam \update_jdo_strobe~0 .lut_mask = 16'hAAFF;
defparam \update_jdo_strobe~0 .sum_lutc_input = "datac";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cycloneive_lcell_comb \jxuir~0 (
	.dataa(\the_altera_std_synchronizer4|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_uir~q ),
	.cin(gnd),
	.combout(\jxuir~0_combout ),
	.cout());
defparam \jxuir~0 .lut_mask = 16'hAAFF;
defparam \jxuir~0 .sum_lutc_input = "datac";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(\ir[1]~q ),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\enable_action_strobe~q ),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(\ir[0]~q ),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_17 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_18 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_debug_slave_tck (
	sr_0,
	MonDReg_0,
	MonDReg_2,
	sr_35,
	MonDReg_3,
	sr_31,
	MonDReg_4,
	MonDReg_29,
	MonDReg_28,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_18,
	MonDReg_10,
	MonDReg_8,
	sr_7,
	sr_15,
	ir_out_0,
	ir_out_1,
	sr_1,
	virtual_state_cdr,
	virtual_state_sdr,
	sr_2,
	break_readreg_0,
	virtual_state_uir,
	hbreak_enabled,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	monitor_ready,
	sr_4,
	break_readreg_2,
	sr_37,
	sr_36,
	sr_17,
	sr_34,
	sr_21,
	sr_20,
	monitor_error,
	sr_5,
	break_readreg_3,
	sr_26,
	sr_28,
	sr_27,
	sr_25,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_19,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_6,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	MonDReg_26,
	break_readreg_24,
	MonDReg_24,
	break_readreg_17,
	MonDReg_17,
	resetlatch,
	break_readreg_31,
	MonDReg_31,
	break_readreg_30,
	MonDReg_30,
	break_readreg_29,
	break_readreg_28,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_21,
	MonDReg_9,
	MonDReg_23,
	MonDReg_22,
	MonDReg_7,
	MonDReg_6,
	break_readreg_18,
	sr_23,
	break_readreg_21,
	break_readreg_5,
	sr_16,
	sr_24,
	break_readreg_22,
	break_readreg_6,
	sr_8,
	break_readreg_15,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_0;
input 	MonDReg_2;
output 	sr_35;
input 	MonDReg_3;
output 	sr_31;
input 	MonDReg_4;
input 	MonDReg_29;
input 	MonDReg_28;
input 	MonDReg_11;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_18;
input 	MonDReg_10;
input 	MonDReg_8;
output 	sr_7;
output 	sr_15;
output 	ir_out_0;
output 	ir_out_1;
output 	sr_1;
input 	virtual_state_cdr;
input 	virtual_state_sdr;
output 	sr_2;
input 	break_readreg_0;
input 	virtual_state_uir;
input 	hbreak_enabled;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
input 	monitor_ready;
output 	sr_4;
input 	break_readreg_2;
output 	sr_37;
output 	sr_36;
output 	sr_17;
output 	sr_34;
output 	sr_21;
output 	sr_20;
input 	monitor_error;
output 	sr_5;
input 	break_readreg_3;
output 	sr_26;
output 	sr_28;
output 	sr_27;
output 	sr_25;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
output 	sr_33;
output 	sr_32;
output 	sr_30;
output 	sr_29;
output 	sr_19;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_17;
input 	MonDReg_17;
input 	resetlatch;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_21;
input 	MonDReg_9;
input 	MonDReg_23;
input 	MonDReg_22;
input 	MonDReg_7;
input 	MonDReg_6;
input 	break_readreg_18;
output 	sr_23;
input 	break_readreg_21;
input 	break_readreg_5;
output 	sr_16;
output 	sr_24;
input 	break_readreg_22;
input 	break_readreg_6;
output 	sr_8;
input 	break_readreg_15;
output 	sr_14;
output 	sr_13;
output 	sr_12;
output 	sr_11;
output 	sr_10;
output 	sr_9;
input 	break_readreg_23;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \DRsize.000~q ;
wire \sr[0]~5_combout ;
wire \Mux37~0_combout ;
wire \sr~10_combout ;
wire \DRsize.100~q ;
wire \sr[35]~6_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr[31]~50_combout ;
wire \sr[31]~7_combout ;
wire \Mux30~0_combout ;
wire \sr[7]~8_combout ;
wire \sr[33]~83_combout ;
wire \DRsize.010~q ;
wire \sr[15]~9_combout ;
wire \sr~71_combout ;
wire \sr~72_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr[5]~13_combout ;
wire \sr~14_combout ;
wire \sr~15_combout ;
wire \sr~16_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr~19_combout ;
wire \sr~20_combout ;
wire \sr[37]~21_combout ;
wire \sr~22_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr[33]~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~55_combout ;
wire \sr~56_combout ;
wire \sr~57_combout ;
wire \sr~58_combout ;
wire \sr~59_combout ;
wire \sr~60_combout ;
wire \sr~61_combout ;
wire \sr~62_combout ;
wire \sr~63_combout ;
wire \sr~64_combout ;
wire \sr~65_combout ;
wire \sr~66_combout ;
wire \sr~67_combout ;
wire \sr~68_combout ;
wire \sr~69_combout ;
wire \sr~70_combout ;
wire \sr~73_combout ;
wire \sr~74_combout ;
wire \sr~75_combout ;
wire \sr~76_combout ;
wire \sr~77_combout ;
wire \sr~78_combout ;
wire \sr~79_combout ;
wire \sr~80_combout ;
wire \sr~81_combout ;
wire \sr~82_combout ;


final_project_soc_altera_std_synchronizer_20 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

final_project_soc_altera_std_synchronizer_19 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr[0]~5_combout ),
	.asdata(\sr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr[35]~6_combout ),
	.asdata(\sr~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr[31]~7_combout ),
	.asdata(sr_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr[7]~8_combout ),
	.asdata(sr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr[15]~9_combout ),
	.asdata(\sr~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[5]~13_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cycloneive_lcell_comb \sr[0]~5 (
	.dataa(altera_internal_jtag1),
	.datab(sr_1),
	.datac(gnd),
	.datad(\DRsize.000~q ),
	.cin(gnd),
	.combout(\sr[0]~5_combout ),
	.cout());
defparam \sr[0]~5 .lut_mask = 16'hAACC;
defparam \sr[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux37~0 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
defparam \Mux37~0 .lut_mask = 16'h7777;
defparam \Mux37~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~10 (
	.dataa(sr_0),
	.datab(virtual_state_cdr),
	.datac(\the_altera_std_synchronizer2|dreg[0]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~10_combout ),
	.cout());
defparam \sr~10 .lut_mask = 16'hFFB8;
defparam \sr~10 .sum_lutc_input = "datac";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cycloneive_lcell_comb \sr[35]~6 (
	.dataa(sr_36),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.100~q ),
	.cin(gnd),
	.combout(\sr[35]~6_combout ),
	.cout());
defparam \sr[35]~6 .lut_mask = 16'hAACC;
defparam \sr[35]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~23 (
	.dataa(irf_reg_1_2),
	.datab(state_3),
	.datac(splitter_nodes_receive_1_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~23_combout ),
	.cout());
defparam \sr~23 .lut_mask = 16'hFDFF;
defparam \sr~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~24 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(sr_35),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr~24_combout ),
	.cout());
defparam \sr~24 .lut_mask = 16'hFFFE;
defparam \sr~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~25 (
	.dataa(irf_reg_0_2),
	.datab(\the_altera_std_synchronizer1|dreg[0]~q ),
	.datac(\sr~23_combout ),
	.datad(\sr~24_combout ),
	.cin(gnd),
	.combout(\sr~25_combout ),
	.cout());
defparam \sr~25 .lut_mask = 16'hFFFD;
defparam \sr~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~50 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(break_readreg_30),
	.datad(MonDReg_30),
	.cin(gnd),
	.combout(\sr[31]~50_combout ),
	.cout());
defparam \sr[31]~50 .lut_mask = 16'hFFF6;
defparam \sr[31]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~7 (
	.dataa(sr_31),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(\sr[31]~50_combout ),
	.cin(gnd),
	.combout(\sr[31]~7_combout ),
	.cout());
defparam \sr[31]~7 .lut_mask = 16'hBF8F;
defparam \sr[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~0 (
	.dataa(break_readreg_6),
	.datab(MonDReg_6),
	.datac(irf_reg_1_2),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hACFF;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[7]~8 (
	.dataa(\Mux30~0_combout ),
	.datab(sr_7),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr[7]~8_combout ),
	.cout());
defparam \sr[7]~8 .lut_mask = 16'hAACC;
defparam \sr[7]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[33]~83 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sr[33]~83_combout ),
	.cout());
defparam \sr[33]~83 .lut_mask = 16'hEEEE;
defparam \sr[33]~83 .sum_lutc_input = "datac";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[33]~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cycloneive_lcell_comb \sr[15]~9 (
	.dataa(sr_16),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.010~q ),
	.cin(gnd),
	.combout(\sr[15]~9_combout ),
	.cout());
defparam \sr[15]~9 .lut_mask = 16'hAACC;
defparam \sr[15]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~71 (
	.dataa(break_readreg_14),
	.datab(MonDReg_14),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~71_combout ),
	.cout());
defparam \sr~71 .lut_mask = 16'hAACC;
defparam \sr~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~72 (
	.dataa(sr_15),
	.datab(virtual_state_cdr),
	.datac(\sr~71_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~72_combout ),
	.cout());
defparam \sr~72 .lut_mask = 16'hB8FF;
defparam \sr~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~11 (
	.dataa(break_readreg_0),
	.datab(MonDReg_0),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~11_combout ),
	.cout());
defparam \sr~11 .lut_mask = 16'hAACC;
defparam \sr~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~12 (
	.dataa(sr_2),
	.datab(virtual_state_sdr),
	.datac(\sr~11_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~12_combout ),
	.cout());
defparam \sr~12 .lut_mask = 16'hB8FF;
defparam \sr~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[5]~13 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr[5]~13_combout ),
	.cout());
defparam \sr[5]~13 .lut_mask = 16'hFEFF;
defparam \sr[5]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~14 (
	.dataa(break_readreg_1),
	.datab(MonDReg_1),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~14_combout ),
	.cout());
defparam \sr~14 .lut_mask = 16'hAACC;
defparam \sr~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~15 (
	.dataa(sr_3),
	.datab(virtual_state_sdr),
	.datac(\sr~14_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~15_combout ),
	.cout());
defparam \sr~15 .lut_mask = 16'hB8FF;
defparam \sr~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~16 (
	.dataa(break_readreg_2),
	.datab(MonDReg_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~16_combout ),
	.cout());
defparam \sr~16 .lut_mask = 16'hAACC;
defparam \sr~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~17 (
	.dataa(sr_4),
	.datab(virtual_state_sdr),
	.datac(\sr~16_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~17_combout ),
	.cout());
defparam \sr~17 .lut_mask = 16'hB8FF;
defparam \sr~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~18 (
	.dataa(break_readreg_3),
	.datab(MonDReg_3),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~18_combout ),
	.cout());
defparam \sr~18 .lut_mask = 16'hAACC;
defparam \sr~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~19 (
	.dataa(sr_5),
	.datab(virtual_state_sdr),
	.datac(\sr~18_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~19_combout ),
	.cout());
defparam \sr~19 .lut_mask = 16'hB8FF;
defparam \sr~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~20 (
	.dataa(altera_internal_jtag1),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~20_combout ),
	.cout());
defparam \sr~20 .lut_mask = 16'hFEFF;
defparam \sr~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[37]~21 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[37]~21_combout ),
	.cout());
defparam \sr[37]~21 .lut_mask = 16'hFF7D;
defparam \sr[37]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~22 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(sr_37),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~22_combout ),
	.cout());
defparam \sr~22 .lut_mask = 16'hFEFF;
defparam \sr~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~26 (
	.dataa(break_readreg_16),
	.datab(MonDReg_16),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~26_combout ),
	.cout());
defparam \sr~26 .lut_mask = 16'hAACC;
defparam \sr~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~27 (
	.dataa(virtual_state_sdr),
	.datab(irf_reg_0_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~27_combout ),
	.cout());
defparam \sr~27 .lut_mask = 16'hEEFF;
defparam \sr~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~28 (
	.dataa(virtual_state_sdr),
	.datab(sr_18),
	.datac(\sr~26_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~28_combout ),
	.cout());
defparam \sr~28 .lut_mask = 16'hFEFF;
defparam \sr~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[33]~29 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[33]~29_combout ),
	.cout());
defparam \sr[33]~29 .lut_mask = 16'hFF7F;
defparam \sr[33]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~30 (
	.dataa(sr_35),
	.datab(virtual_state_sdr),
	.datac(monitor_error),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~30_combout ),
	.cout());
defparam \sr~30 .lut_mask = 16'hFFB8;
defparam \sr~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~31 (
	.dataa(break_readreg_20),
	.datab(MonDReg_20),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~31_combout ),
	.cout());
defparam \sr~31 .lut_mask = 16'hAACC;
defparam \sr~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~32 (
	.dataa(virtual_state_sdr),
	.datab(sr_22),
	.datac(\sr~31_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~32_combout ),
	.cout());
defparam \sr~32 .lut_mask = 16'hFEFF;
defparam \sr~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~33 (
	.dataa(break_readreg_19),
	.datab(MonDReg_19),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~33_combout ),
	.cout());
defparam \sr~33 .lut_mask = 16'hAACC;
defparam \sr~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~34 (
	.dataa(virtual_state_sdr),
	.datab(sr_21),
	.datac(\sr~33_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~34_combout ),
	.cout());
defparam \sr~34 .lut_mask = 16'hFEFF;
defparam \sr~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~35 (
	.dataa(break_readreg_4),
	.datab(MonDReg_4),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~35_combout ),
	.cout());
defparam \sr~35 .lut_mask = 16'hAACC;
defparam \sr~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~36 (
	.dataa(sr_6),
	.datab(virtual_state_sdr),
	.datac(\sr~35_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~36_combout ),
	.cout());
defparam \sr~36 .lut_mask = 16'hB8FF;
defparam \sr~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~37 (
	.dataa(break_readreg_25),
	.datab(MonDReg_25),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~37_combout ),
	.cout());
defparam \sr~37 .lut_mask = 16'hAACC;
defparam \sr~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~38 (
	.dataa(virtual_state_sdr),
	.datab(sr_27),
	.datac(\sr~37_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~38_combout ),
	.cout());
defparam \sr~38 .lut_mask = 16'hFEFF;
defparam \sr~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~39 (
	.dataa(break_readreg_27),
	.datab(MonDReg_27),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~39_combout ),
	.cout());
defparam \sr~39 .lut_mask = 16'hAACC;
defparam \sr~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~40 (
	.dataa(virtual_state_sdr),
	.datab(sr_29),
	.datac(\sr~39_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~40_combout ),
	.cout());
defparam \sr~40 .lut_mask = 16'hFEFF;
defparam \sr~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~41 (
	.dataa(break_readreg_26),
	.datab(MonDReg_26),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~41_combout ),
	.cout());
defparam \sr~41 .lut_mask = 16'hAACC;
defparam \sr~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~42 (
	.dataa(virtual_state_sdr),
	.datab(sr_28),
	.datac(\sr~41_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~42_combout ),
	.cout());
defparam \sr~42 .lut_mask = 16'hFEFF;
defparam \sr~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~43 (
	.dataa(break_readreg_24),
	.datab(MonDReg_24),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~43_combout ),
	.cout());
defparam \sr~43 .lut_mask = 16'hAACC;
defparam \sr~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~44 (
	.dataa(virtual_state_sdr),
	.datab(sr_26),
	.datac(\sr~43_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~44_combout ),
	.cout());
defparam \sr~44 .lut_mask = 16'hFEFF;
defparam \sr~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~45 (
	.dataa(break_readreg_17),
	.datab(MonDReg_17),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~45_combout ),
	.cout());
defparam \sr~45 .lut_mask = 16'hAACC;
defparam \sr~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~46 (
	.dataa(virtual_state_sdr),
	.datab(sr_19),
	.datac(\sr~45_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~46_combout ),
	.cout());
defparam \sr~46 .lut_mask = 16'hFEFF;
defparam \sr~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~47 (
	.dataa(sr_34),
	.datab(virtual_state_sdr),
	.datac(resetlatch),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~47_combout ),
	.cout());
defparam \sr~47 .lut_mask = 16'hFFB8;
defparam \sr~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~48 (
	.dataa(break_readreg_31),
	.datab(MonDReg_31),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~48_combout ),
	.cout());
defparam \sr~48 .lut_mask = 16'hAACC;
defparam \sr~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~49 (
	.dataa(virtual_state_sdr),
	.datab(sr_33),
	.datac(\sr~48_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~49_combout ),
	.cout());
defparam \sr~49 .lut_mask = 16'hFEFF;
defparam \sr~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~51 (
	.dataa(break_readreg_29),
	.datab(MonDReg_29),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~51_combout ),
	.cout());
defparam \sr~51 .lut_mask = 16'hAACC;
defparam \sr~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~52 (
	.dataa(virtual_state_sdr),
	.datab(sr_31),
	.datac(\sr~51_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~52_combout ),
	.cout());
defparam \sr~52 .lut_mask = 16'hFEFF;
defparam \sr~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~53 (
	.dataa(break_readreg_28),
	.datab(MonDReg_28),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~53_combout ),
	.cout());
defparam \sr~53 .lut_mask = 16'hAACC;
defparam \sr~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~54 (
	.dataa(virtual_state_sdr),
	.datab(sr_30),
	.datac(\sr~53_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~54_combout ),
	.cout());
defparam \sr~54 .lut_mask = 16'hFEFF;
defparam \sr~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~55 (
	.dataa(break_readreg_18),
	.datab(MonDReg_18),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~55_combout ),
	.cout());
defparam \sr~55 .lut_mask = 16'hAACC;
defparam \sr~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~56 (
	.dataa(virtual_state_sdr),
	.datab(sr_20),
	.datac(\sr~55_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~56_combout ),
	.cout());
defparam \sr~56 .lut_mask = 16'hFEFF;
defparam \sr~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~57 (
	.dataa(break_readreg_21),
	.datab(MonDReg_21),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~57_combout ),
	.cout());
defparam \sr~57 .lut_mask = 16'hAACC;
defparam \sr~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~58 (
	.dataa(virtual_state_sdr),
	.datab(sr_23),
	.datac(\sr~57_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~58_combout ),
	.cout());
defparam \sr~58 .lut_mask = 16'hFEFF;
defparam \sr~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~59 (
	.dataa(break_readreg_5),
	.datab(MonDReg_5),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~59_combout ),
	.cout());
defparam \sr~59 .lut_mask = 16'hAACC;
defparam \sr~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~60 (
	.dataa(sr_7),
	.datab(virtual_state_sdr),
	.datac(\sr~59_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~60_combout ),
	.cout());
defparam \sr~60 .lut_mask = 16'hB8FF;
defparam \sr~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~61 (
	.dataa(break_readreg_22),
	.datab(MonDReg_22),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~61_combout ),
	.cout());
defparam \sr~61 .lut_mask = 16'hAACC;
defparam \sr~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~62 (
	.dataa(virtual_state_sdr),
	.datab(sr_24),
	.datac(\sr~61_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~62_combout ),
	.cout());
defparam \sr~62 .lut_mask = 16'hFEFF;
defparam \sr~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~63 (
	.dataa(break_readreg_15),
	.datab(MonDReg_15),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~63_combout ),
	.cout());
defparam \sr~63 .lut_mask = 16'hAACC;
defparam \sr~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~64 (
	.dataa(virtual_state_sdr),
	.datab(sr_17),
	.datac(\sr~63_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~64_combout ),
	.cout());
defparam \sr~64 .lut_mask = 16'hFEFF;
defparam \sr~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~65 (
	.dataa(break_readreg_23),
	.datab(MonDReg_23),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~65_combout ),
	.cout());
defparam \sr~65 .lut_mask = 16'hAACC;
defparam \sr~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~66 (
	.dataa(virtual_state_sdr),
	.datab(sr_25),
	.datac(\sr~65_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~66_combout ),
	.cout());
defparam \sr~66 .lut_mask = 16'hFEFF;
defparam \sr~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~67 (
	.dataa(break_readreg_7),
	.datab(MonDReg_7),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~67_combout ),
	.cout());
defparam \sr~67 .lut_mask = 16'hAACC;
defparam \sr~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~68 (
	.dataa(sr_9),
	.datab(virtual_state_sdr),
	.datac(\sr~67_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~68_combout ),
	.cout());
defparam \sr~68 .lut_mask = 16'hB8FF;
defparam \sr~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~69 (
	.dataa(break_readreg_13),
	.datab(MonDReg_13),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~69_combout ),
	.cout());
defparam \sr~69 .lut_mask = 16'hAACC;
defparam \sr~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~70 (
	.dataa(sr_15),
	.datab(virtual_state_sdr),
	.datac(\sr~69_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~70_combout ),
	.cout());
defparam \sr~70 .lut_mask = 16'hB8FF;
defparam \sr~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~73 (
	.dataa(break_readreg_12),
	.datab(MonDReg_12),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~73_combout ),
	.cout());
defparam \sr~73 .lut_mask = 16'hAACC;
defparam \sr~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~74 (
	.dataa(sr_14),
	.datab(virtual_state_sdr),
	.datac(\sr~73_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~74_combout ),
	.cout());
defparam \sr~74 .lut_mask = 16'hB8FF;
defparam \sr~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~75 (
	.dataa(break_readreg_11),
	.datab(MonDReg_11),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~75_combout ),
	.cout());
defparam \sr~75 .lut_mask = 16'hAACC;
defparam \sr~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~76 (
	.dataa(sr_13),
	.datab(virtual_state_sdr),
	.datac(\sr~75_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~76_combout ),
	.cout());
defparam \sr~76 .lut_mask = 16'hB8FF;
defparam \sr~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~77 (
	.dataa(break_readreg_10),
	.datab(MonDReg_10),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~77_combout ),
	.cout());
defparam \sr~77 .lut_mask = 16'hAACC;
defparam \sr~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~78 (
	.dataa(sr_12),
	.datab(virtual_state_sdr),
	.datac(\sr~77_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~78_combout ),
	.cout());
defparam \sr~78 .lut_mask = 16'hB8FF;
defparam \sr~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~79 (
	.dataa(break_readreg_9),
	.datab(MonDReg_9),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~79_combout ),
	.cout());
defparam \sr~79 .lut_mask = 16'hAACC;
defparam \sr~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~80 (
	.dataa(sr_11),
	.datab(virtual_state_sdr),
	.datac(\sr~79_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~80_combout ),
	.cout());
defparam \sr~80 .lut_mask = 16'hB8FF;
defparam \sr~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~81 (
	.dataa(break_readreg_8),
	.datab(MonDReg_8),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~81_combout ),
	.cout());
defparam \sr~81 .lut_mask = 16'hAACC;
defparam \sr~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~82 (
	.dataa(sr_10),
	.datab(virtual_state_sdr),
	.datac(\sr~81_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~82_combout ),
	.cout());
defparam \sr~82 .lut_mask = 16'hB8FF;
defparam \sr~82 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_std_synchronizer_19 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_altera_std_synchronizer_20 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_sld_virtual_jtag_basic_1 (
	virtual_state_cdr1,
	virtual_state_sdr,
	virtual_state_uir,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_cdr1;
output 	virtual_state_sdr;
output 	virtual_state_uir;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb virtual_state_cdr(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_3),
	.datad(splitter_nodes_receive_1_3),
	.cin(gnd),
	.combout(virtual_state_cdr1),
	.cout());
defparam virtual_state_cdr.lut_mask = 16'hAFFF;
defparam virtual_state_cdr.sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_sdr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_sdr),
	.cout());
defparam \virtual_state_sdr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_sdr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_uir~0 (
	.dataa(virtual_ir_scan_reg),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(virtual_state_uir),
	.cout());
defparam \virtual_state_uir~0 .lut_mask = 16'hFEFE;
defparam \virtual_state_uir~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_udr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_udr),
	.cout());
defparam \virtual_state_udr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_udr~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	oci_ienable_1,
	oci_ienable_0,
	oci_single_step_mode1,
	debugaccess,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	Equal0,
	take_action_ocireg,
	writedata_1,
	Equal1,
	writedata_3,
	oci_ienable_16,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
output 	oci_ienable_1;
output 	oci_ienable_0;
output 	oci_single_step_mode1;
input 	debugaccess;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
output 	Equal0;
output 	take_action_ocireg;
input 	writedata_1;
output 	Equal1;
input 	writedata_3;
output 	oci_ienable_16;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \oci_ienable[1]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[0]~1_combout ;
wire \oci_single_step_mode~0_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;


dffeas \oci_ienable[1] (
	.clk(clk_clk),
	.d(\oci_ienable[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_1),
	.prn(vcc));
defparam \oci_ienable[1] .is_wysiwyg = "true";
defparam \oci_ienable[1] .power_up = "low";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(\oci_ienable[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(address_0),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocireg~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(Equal0),
	.datad(gnd),
	.cin(gnd),
	.combout(take_action_ocireg),
	.cout());
defparam \take_action_ocireg~0 .lut_mask = 16'hFEFE;
defparam \take_action_ocireg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(address_0),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFE;
defparam \Equal1~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[16] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_16),
	.prn(vcc));
defparam \oci_ienable[16] .is_wysiwyg = "true";
defparam \oci_ienable[16] .power_up = "low";

cycloneive_lcell_comb \oci_ienable[1]~0 (
	.dataa(writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[1]~0_combout ),
	.cout());
defparam \oci_ienable[1]~0 .lut_mask = 16'h5555;
defparam \oci_ienable[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(Equal1),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.cout());
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 16'hFEFE;
defparam \take_action_oci_intr_mask_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[0]~1 (
	.dataa(writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[0]~1_combout ),
	.cout());
defparam \oci_ienable[0]~1 .lut_mask = 16'h5555;
defparam \oci_ienable[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_single_step_mode~0 (
	.dataa(writedata_3),
	.datab(oci_single_step_mode1),
	.datac(gnd),
	.datad(take_action_ocireg),
	.cin(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.cout());
defparam \oci_single_step_mode~0 .lut_mask = 16'hAACC;
defparam \oci_single_step_mode~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(address_8),
	.datab(address_5),
	.datac(address_6),
	.datad(address_7),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hBFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(address_1),
	.datab(address_2),
	.datac(address_3),
	.datad(address_4),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	jdo_0,
	jdo_37,
	jdo_36,
	take_no_action_break_a,
	jdo_3,
	jdo_17,
	jdo_21,
	jdo_20,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_25,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_19,
	jdo_18,
	break_readreg_3,
	jdo_2,
	jdo_5,
	break_readreg_16,
	break_readreg_20,
	break_readreg_19,
	jdo_23,
	break_readreg_4,
	jdo_6,
	break_readreg_25,
	break_readreg_27,
	break_readreg_26,
	break_readreg_24,
	break_readreg_17,
	jdo_16,
	break_readreg_31,
	break_readreg_30,
	break_readreg_29,
	break_readreg_28,
	break_readreg_18,
	break_readreg_21,
	jdo_22,
	jdo_7,
	break_readreg_5,
	jdo_24,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_22,
	break_readreg_6,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
input 	jdo_0;
input 	jdo_37;
input 	jdo_36;
input 	take_no_action_break_a;
input 	jdo_3;
input 	jdo_17;
input 	jdo_21;
input 	jdo_20;
output 	break_readreg_2;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_25;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
input 	jdo_19;
input 	jdo_18;
output 	break_readreg_3;
input 	jdo_2;
input 	jdo_5;
output 	break_readreg_16;
output 	break_readreg_20;
output 	break_readreg_19;
input 	jdo_23;
output 	break_readreg_4;
input 	jdo_6;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_24;
output 	break_readreg_17;
input 	jdo_16;
output 	break_readreg_31;
output 	break_readreg_30;
output 	break_readreg_29;
output 	break_readreg_28;
output 	break_readreg_18;
output 	break_readreg_21;
input 	jdo_22;
input 	jdo_7;
output 	break_readreg_5;
input 	jdo_24;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
output 	break_readreg_22;
output 	break_readreg_6;
output 	break_readreg_15;
output 	break_readreg_23;
output 	break_readreg_7;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_10;
output 	break_readreg_9;
output 	break_readreg_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg~0_combout ;
wire \break_readreg~1_combout ;
wire \break_readreg~2_combout ;
wire \break_readreg~3_combout ;
wire \break_readreg~4_combout ;
wire \break_readreg~5_combout ;
wire \break_readreg~6_combout ;
wire \break_readreg~7_combout ;
wire \break_readreg~8_combout ;
wire \break_readreg~9_combout ;
wire \break_readreg~10_combout ;
wire \break_readreg~11_combout ;
wire \break_readreg~12_combout ;
wire \break_readreg~13_combout ;
wire \break_readreg~14_combout ;
wire \break_readreg~15_combout ;
wire \break_readreg~16_combout ;
wire \break_readreg~17_combout ;
wire \break_readreg~18_combout ;
wire \break_readreg~19_combout ;
wire \break_readreg~20_combout ;
wire \break_readreg~21_combout ;
wire \break_readreg~22_combout ;
wire \break_readreg~23_combout ;
wire \break_readreg~24_combout ;
wire \break_readreg~25_combout ;
wire \break_readreg~26_combout ;
wire \break_readreg~27_combout ;
wire \break_readreg~28_combout ;
wire \break_readreg~29_combout ;
wire \break_readreg~30_combout ;
wire \break_readreg~31_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(\break_readreg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(\break_readreg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(\break_readreg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(\break_readreg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(\break_readreg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(\break_readreg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(\break_readreg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(\break_readreg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(\break_readreg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(\break_readreg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(\break_readreg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(\break_readreg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(\break_readreg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(\break_readreg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(\break_readreg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(\break_readreg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(\break_readreg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(\break_readreg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(\break_readreg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(\break_readreg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(\break_readreg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(\break_readreg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(\break_readreg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(\break_readreg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(\break_readreg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(\break_readreg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(\break_readreg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(\break_readreg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(\break_readreg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(\break_readreg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(\break_readreg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(\break_readreg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_no_action_break_a),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

cycloneive_lcell_comb \break_readreg~0 (
	.dataa(jdo_0),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~0_combout ),
	.cout());
defparam \break_readreg~0 .lut_mask = 16'hFEFF;
defparam \break_readreg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~1 (
	.dataa(jdo_1),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~1_combout ),
	.cout());
defparam \break_readreg~1 .lut_mask = 16'hFEFF;
defparam \break_readreg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~2 (
	.dataa(jdo_2),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~2_combout ),
	.cout());
defparam \break_readreg~2 .lut_mask = 16'hFEFF;
defparam \break_readreg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~3 (
	.dataa(jdo_3),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~3_combout ),
	.cout());
defparam \break_readreg~3 .lut_mask = 16'hFEFF;
defparam \break_readreg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~4 (
	.dataa(jdo_16),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~4_combout ),
	.cout());
defparam \break_readreg~4 .lut_mask = 16'hFEFF;
defparam \break_readreg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~5 (
	.dataa(jdo_20),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~5_combout ),
	.cout());
defparam \break_readreg~5 .lut_mask = 16'hFEFF;
defparam \break_readreg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~6 (
	.dataa(jdo_19),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~6_combout ),
	.cout());
defparam \break_readreg~6 .lut_mask = 16'hFEFF;
defparam \break_readreg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~7 (
	.dataa(jdo_4),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~7_combout ),
	.cout());
defparam \break_readreg~7 .lut_mask = 16'hFEFF;
defparam \break_readreg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~8 (
	.dataa(jdo_25),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~8_combout ),
	.cout());
defparam \break_readreg~8 .lut_mask = 16'hFEFF;
defparam \break_readreg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~9 (
	.dataa(jdo_27),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~9_combout ),
	.cout());
defparam \break_readreg~9 .lut_mask = 16'hFEFF;
defparam \break_readreg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~10 (
	.dataa(jdo_26),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~10_combout ),
	.cout());
defparam \break_readreg~10 .lut_mask = 16'hFEFF;
defparam \break_readreg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~11 (
	.dataa(jdo_24),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~11_combout ),
	.cout());
defparam \break_readreg~11 .lut_mask = 16'hFEFF;
defparam \break_readreg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~12 (
	.dataa(jdo_17),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~12_combout ),
	.cout());
defparam \break_readreg~12 .lut_mask = 16'hFEFF;
defparam \break_readreg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~13 (
	.dataa(jdo_31),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~13_combout ),
	.cout());
defparam \break_readreg~13 .lut_mask = 16'hFEFF;
defparam \break_readreg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~14 (
	.dataa(jdo_30),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~14_combout ),
	.cout());
defparam \break_readreg~14 .lut_mask = 16'hFEFF;
defparam \break_readreg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~15 (
	.dataa(jdo_29),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~15_combout ),
	.cout());
defparam \break_readreg~15 .lut_mask = 16'hFEFF;
defparam \break_readreg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~16 (
	.dataa(jdo_28),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~16_combout ),
	.cout());
defparam \break_readreg~16 .lut_mask = 16'hFEFF;
defparam \break_readreg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~17 (
	.dataa(jdo_18),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~17_combout ),
	.cout());
defparam \break_readreg~17 .lut_mask = 16'hFEFF;
defparam \break_readreg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~18 (
	.dataa(jdo_21),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~18_combout ),
	.cout());
defparam \break_readreg~18 .lut_mask = 16'hFEFF;
defparam \break_readreg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~19 (
	.dataa(jdo_5),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~19_combout ),
	.cout());
defparam \break_readreg~19 .lut_mask = 16'hFEFF;
defparam \break_readreg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~20 (
	.dataa(jdo_22),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~20_combout ),
	.cout());
defparam \break_readreg~20 .lut_mask = 16'hFEFF;
defparam \break_readreg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~21 (
	.dataa(jdo_6),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~21_combout ),
	.cout());
defparam \break_readreg~21 .lut_mask = 16'hFEFF;
defparam \break_readreg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~22 (
	.dataa(jdo_15),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~22_combout ),
	.cout());
defparam \break_readreg~22 .lut_mask = 16'hFEFF;
defparam \break_readreg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~23 (
	.dataa(jdo_23),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~23_combout ),
	.cout());
defparam \break_readreg~23 .lut_mask = 16'hFEFF;
defparam \break_readreg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~24 (
	.dataa(jdo_7),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~24_combout ),
	.cout());
defparam \break_readreg~24 .lut_mask = 16'hFEFF;
defparam \break_readreg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~25 (
	.dataa(jdo_13),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~25_combout ),
	.cout());
defparam \break_readreg~25 .lut_mask = 16'hFEFF;
defparam \break_readreg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~26 (
	.dataa(jdo_14),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~26_combout ),
	.cout());
defparam \break_readreg~26 .lut_mask = 16'hFEFF;
defparam \break_readreg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~27 (
	.dataa(jdo_12),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~27_combout ),
	.cout());
defparam \break_readreg~27 .lut_mask = 16'hFEFF;
defparam \break_readreg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~28 (
	.dataa(jdo_11),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~28_combout ),
	.cout());
defparam \break_readreg~28 .lut_mask = 16'hFEFF;
defparam \break_readreg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~29 (
	.dataa(jdo_10),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~29_combout ),
	.cout());
defparam \break_readreg~29 .lut_mask = 16'hFEFF;
defparam \break_readreg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~30 (
	.dataa(jdo_9),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~30_combout ),
	.cout());
defparam \break_readreg~30 .lut_mask = 16'hFEFF;
defparam \break_readreg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~31 (
	.dataa(jdo_8),
	.datab(jdo_37),
	.datac(jdo_36),
	.datad(take_no_action_break_a),
	.cin(gnd),
	.combout(\break_readreg~31_combout ),
	.cout());
defparam \break_readreg~31 .lut_mask = 16'hFEFF;
defparam \break_readreg~31 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_oci_debug (
	jtag_break1,
	r_sync_rst,
	jdo_35,
	take_action_ocimem_a,
	monitor_ready1,
	jdo_34,
	jdo_21,
	jdo_20,
	take_action_ocimem_a1,
	writedata_0,
	take_action_ocireg,
	jdo_25,
	writedata_1,
	jdo_19,
	jdo_18,
	monitor_error1,
	monitor_go1,
	jdo_23,
	resetlatch1,
	jdo_24,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	jtag_break1;
input 	r_sync_rst;
input 	jdo_35;
input 	take_action_ocimem_a;
output 	monitor_ready1;
input 	jdo_34;
input 	jdo_21;
input 	jdo_20;
input 	take_action_ocimem_a1;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_25;
input 	writedata_1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_error1;
output 	monitor_go1;
input 	jdo_23;
output 	resetlatch1;
input 	jdo_24;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \jtag_break~1_combout ;
wire \always1~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


final_project_soc_altera_std_synchronizer_21 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(\jtag_break~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cycloneive_lcell_comb \break_on_reset~0 (
	.dataa(\break_on_reset~q ),
	.datab(jdo_19),
	.datac(jdo_18),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\break_on_reset~0_combout ),
	.cout());
defparam \break_on_reset~0 .lut_mask = 16'hAFCF;
defparam \break_on_reset~0 .sum_lutc_input = "datac";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cycloneive_lcell_comb \jtag_break~0 (
	.dataa(jtag_break1),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(\the_altera_std_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\jtag_break~0_combout ),
	.cout());
defparam \jtag_break~0 .lut_mask = 16'hAACC;
defparam \jtag_break~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_break~1 (
	.dataa(jdo_21),
	.datab(jtag_break1),
	.datac(gnd),
	.datad(jdo_20),
	.cin(gnd),
	.combout(\jtag_break~1_combout ),
	.cout());
defparam \jtag_break~1 .lut_mask = 16'hEEFF;
defparam \jtag_break~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(take_action_ocimem_a),
	.datab(jdo_34),
	.datac(jdo_25),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFF;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_ready~0 (
	.dataa(monitor_ready1),
	.datab(writedata_0),
	.datac(take_action_ocireg),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_ready~0_combout ),
	.cout());
defparam \monitor_ready~0 .lut_mask = 16'hFEFF;
defparam \monitor_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_error~0 (
	.dataa(monitor_error1),
	.datab(take_action_ocireg),
	.datac(writedata_1),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_error~0_combout ),
	.cout());
defparam \monitor_error~0 .lut_mask = 16'hFEFF;
defparam \monitor_error~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_go~0 (
	.dataa(jdo_23),
	.datab(monitor_go1),
	.datac(take_action_ocimem_a1),
	.datad(state_1),
	.cin(gnd),
	.combout(\monitor_go~0_combout ),
	.cout());
defparam \monitor_go~0 .lut_mask = 16'hFEFF;
defparam \monitor_go~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \resetlatch~0 (
	.dataa(take_action_ocimem_a1),
	.datab(resetlatch1),
	.datac(\the_altera_std_synchronizer|dreg[0]~q ),
	.datad(jdo_24),
	.cin(gnd),
	.combout(\resetlatch~0_combout ),
	.cout());
defparam \resetlatch~0 .lut_mask = 16'hFDFF;
defparam \resetlatch~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altera_std_synchronizer_21 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem (
	MonDReg_0,
	q_a_0,
	MonDReg_2,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	MonDReg_3,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_31,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_10,
	q_a_24,
	q_a_9,
	q_a_23,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	MonDReg_4,
	MonDReg_29,
	MonDReg_28,
	MonDReg_11,
	MonDReg_12,
	MonDReg_5,
	MonDReg_18,
	MonDReg_10,
	MonDReg_8,
	waitrequest1,
	write,
	address_8,
	read,
	MonDReg_1,
	jdo_3,
	jdo_35,
	take_action_ocimem_b,
	take_action_ocimem_a,
	jdo_17,
	jdo_34,
	jdo_21,
	jdo_20,
	take_action_ocimem_a1,
	r_early_rst,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	debugaccess,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	byteenable_0,
	jdo_25,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	writedata_1,
	jdo_19,
	jdo_18,
	writedata_3,
	jdo_5,
	MonDReg_16,
	MonDReg_20,
	MonDReg_19,
	jdo_23,
	writedata_2,
	writedata_4,
	jdo_6,
	MonDReg_25,
	MonDReg_27,
	MonDReg_26,
	MonDReg_24,
	MonDReg_17,
	jdo_16,
	MonDReg_31,
	MonDReg_30,
	writedata_11,
	byteenable_1,
	MonDReg_13,
	writedata_13,
	writedata_16,
	byteenable_2,
	writedata_12,
	writedata_5,
	MonDReg_14,
	writedata_14,
	MonDReg_15,
	writedata_15,
	MonDReg_21,
	writedata_21,
	writedata_18,
	writedata_17,
	writedata_31,
	byteenable_3,
	writedata_30,
	writedata_29,
	writedata_28,
	writedata_27,
	writedata_26,
	writedata_25,
	writedata_10,
	writedata_24,
	MonDReg_9,
	writedata_9,
	MonDReg_23,
	writedata_23,
	writedata_8,
	MonDReg_22,
	writedata_22,
	MonDReg_7,
	writedata_7,
	MonDReg_6,
	writedata_6,
	writedata_20,
	writedata_19,
	jdo_22,
	jdo_7,
	jdo_24,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_0;
output 	q_a_0;
output 	MonDReg_2;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	MonDReg_3;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_31;
output 	q_a_30;
output 	q_a_29;
output 	q_a_28;
output 	q_a_27;
output 	q_a_26;
output 	q_a_25;
output 	q_a_10;
output 	q_a_24;
output 	q_a_9;
output 	q_a_23;
output 	q_a_8;
output 	q_a_22;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_19;
output 	MonDReg_4;
output 	MonDReg_29;
output 	MonDReg_28;
output 	MonDReg_11;
output 	MonDReg_12;
output 	MonDReg_5;
output 	MonDReg_18;
output 	MonDReg_10;
output 	MonDReg_8;
output 	waitrequest1;
input 	write;
input 	address_8;
input 	read;
output 	MonDReg_1;
input 	jdo_3;
input 	jdo_35;
input 	take_action_ocimem_b;
input 	take_action_ocimem_a;
input 	jdo_17;
input 	jdo_34;
input 	jdo_21;
input 	jdo_20;
input 	take_action_ocimem_a1;
input 	r_early_rst;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	debugaccess;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
input 	byteenable_0;
input 	jdo_25;
input 	jdo_33;
input 	jdo_32;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
input 	writedata_1;
input 	jdo_19;
input 	jdo_18;
input 	writedata_3;
input 	jdo_5;
output 	MonDReg_16;
output 	MonDReg_20;
output 	MonDReg_19;
input 	jdo_23;
input 	writedata_2;
input 	writedata_4;
input 	jdo_6;
output 	MonDReg_25;
output 	MonDReg_27;
output 	MonDReg_26;
output 	MonDReg_24;
output 	MonDReg_17;
input 	jdo_16;
output 	MonDReg_31;
output 	MonDReg_30;
input 	writedata_11;
input 	byteenable_1;
output 	MonDReg_13;
input 	writedata_13;
input 	writedata_16;
input 	byteenable_2;
input 	writedata_12;
input 	writedata_5;
output 	MonDReg_14;
input 	writedata_14;
output 	MonDReg_15;
input 	writedata_15;
output 	MonDReg_21;
input 	writedata_21;
input 	writedata_18;
input 	writedata_17;
input 	writedata_31;
input 	byteenable_3;
input 	writedata_30;
input 	writedata_29;
input 	writedata_28;
input 	writedata_27;
input 	writedata_26;
input 	writedata_25;
input 	writedata_10;
input 	writedata_24;
output 	MonDReg_9;
input 	writedata_9;
output 	MonDReg_23;
input 	writedata_23;
input 	writedata_8;
output 	MonDReg_22;
input 	writedata_22;
output 	MonDReg_7;
input 	writedata_7;
output 	MonDReg_6;
input 	writedata_6;
input 	writedata_20;
input 	writedata_19;
input 	jdo_22;
input 	jdo_7;
input 	jdo_24;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ociram_wr_en~0_combout ;
wire \jtag_ram_wr~q ;
wire \ociram_wr_en~1_combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[3]~3_combout ;
wire \ociram_wr_data[4]~4_combout ;
wire \ociram_wr_data[11]~5_combout ;
wire \ociram_byteenable[1]~1_combout ;
wire \ociram_wr_data[13]~6_combout ;
wire \ociram_wr_data[16]~7_combout ;
wire \ociram_byteenable[2]~2_combout ;
wire \ociram_wr_data[12]~8_combout ;
wire \ociram_wr_data[5]~9_combout ;
wire \ociram_wr_data[14]~10_combout ;
wire \ociram_wr_data[15]~11_combout ;
wire \ociram_wr_data[21]~12_combout ;
wire \ociram_wr_data[18]~13_combout ;
wire \ociram_wr_data[17]~14_combout ;
wire \ociram_wr_data[31]~15_combout ;
wire \ociram_byteenable[3]~3_combout ;
wire \ociram_wr_data[30]~16_combout ;
wire \ociram_wr_data[29]~17_combout ;
wire \ociram_wr_data[28]~18_combout ;
wire \ociram_wr_data[27]~19_combout ;
wire \ociram_wr_data[26]~20_combout ;
wire \ociram_wr_data[25]~21_combout ;
wire \ociram_wr_data[10]~22_combout ;
wire \ociram_wr_data[24]~23_combout ;
wire \ociram_wr_data[9]~24_combout ;
wire \ociram_wr_data[23]~25_combout ;
wire \ociram_wr_data[8]~26_combout ;
wire \ociram_wr_data[22]~27_combout ;
wire \ociram_wr_data[7]~28_combout ;
wire \ociram_wr_data[6]~29_combout ;
wire \ociram_wr_data[20]~30_combout ;
wire \ociram_wr_data[19]~31_combout ;
wire \MonARegAddrInc[0]~0_combout ;
wire \MonAReg~0_combout ;
wire \MonAReg[2]~q ;
wire \MonARegAddrInc[0]~1 ;
wire \MonARegAddrInc[1]~2_combout ;
wire \MonAReg~2_combout ;
wire \MonAReg[3]~q ;
wire \MonARegAddrInc[1]~3 ;
wire \MonARegAddrInc[2]~4_combout ;
wire \MonAReg~1_combout ;
wire \MonAReg[4]~q ;
wire \Equal0~0_combout ;
wire \MonAReg~3_combout ;
wire \MonAReg[10]~q ;
wire \MonARegAddrInc[2]~5 ;
wire \MonARegAddrInc[3]~6_combout ;
wire \MonAReg~8_combout ;
wire \MonAReg[5]~q ;
wire \MonARegAddrInc[3]~7 ;
wire \MonARegAddrInc[4]~8_combout ;
wire \MonAReg~7_combout ;
wire \MonAReg[6]~q ;
wire \MonARegAddrInc[4]~9 ;
wire \MonARegAddrInc[5]~10_combout ;
wire \MonAReg~6_combout ;
wire \MonAReg[7]~q ;
wire \MonARegAddrInc[5]~11 ;
wire \MonARegAddrInc[6]~12_combout ;
wire \MonAReg~5_combout ;
wire \MonAReg[8]~q ;
wire \MonARegAddrInc[6]~13 ;
wire \MonARegAddrInc[7]~14_combout ;
wire \MonAReg~4_combout ;
wire \MonAReg[9]~q ;
wire \MonARegAddrInc[7]~15 ;
wire \MonARegAddrInc[8]~16_combout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~1_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[0]~0_combout ;
wire \jtag_rd~0_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~12_combout ;
wire \MonDReg[2]~1_combout ;
wire \MonDReg[3]~2_combout ;
wire \MonDReg[4]~3_combout ;
wire \Equal0~1_combout ;
wire \MonDReg[29]~8_combout ;
wire \cfgrom_readdata[28]~0_combout ;
wire \MonDReg[28]~9_combout ;
wire \MonDReg[28]~24_combout ;
wire \MonDReg[11]~5_combout ;
wire \MonDReg[12]~6_combout ;
wire \Equal0~2_combout ;
wire \MonDReg[5]~4_combout ;
wire \Equal0~3_combout ;
wire \MonDReg[18]~7_combout ;
wire \MonDReg[10]~10_combout ;
wire \cfgrom_readdata[8]~1_combout ;
wire \MonDReg[8]~11_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~1_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~1_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~20_combout ;
wire \MonDReg~21_combout ;
wire \MonDReg~22_combout ;
wire \MonDReg~23_combout ;
wire \MonDReg~25_combout ;
wire \MonDReg~26_combout ;
wire \MonDReg~27_combout ;
wire \MonDReg~28_combout ;
wire \MonDReg~29_combout ;
wire \MonDReg~30_combout ;
wire \MonDReg~31_combout ;
wire \MonDReg~32_combout ;
wire \MonDReg~33_combout ;


final_project_soc_final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_5(q_a_5),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_31(q_a_31),
	.q_a_30(q_a_30),
	.q_a_29(q_a_29),
	.q_a_28(q_a_28),
	.q_a_27(q_a_27),
	.q_a_26(q_a_26),
	.q_a_25(q_a_25),
	.q_a_10(q_a_10),
	.q_a_24(q_a_24),
	.q_a_9(q_a_9),
	.q_a_23(q_a_23),
	.q_a_8(q_a_8),
	.q_a_22(q_a_22),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.r_early_rst(r_early_rst),
	.ociram_wr_en(\ociram_wr_en~1_combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~3_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~4_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~5_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~1_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~6_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~7_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~2_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~8_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~9_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~10_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~11_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~12_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~13_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~14_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~15_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~3_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~16_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~17_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~18_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~19_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~20_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~21_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~22_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~23_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~24_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~25_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~26_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~27_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~28_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~29_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~30_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~31_combout ),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \ociram_wr_en~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(address_8),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.cout());
defparam \ociram_wr_en~0 .lut_mask = 16'hEFFF;
defparam \ociram_wr_en~0 .sum_lutc_input = "datac";

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cycloneive_lcell_comb \ociram_wr_en~1 (
	.dataa(\ociram_wr_en~0_combout ),
	.datab(\jtag_ram_access~q ),
	.datac(\jtag_ram_wr~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_wr_en~1_combout ),
	.cout());
defparam \ociram_wr_en~1 .lut_mask = 16'hFEFE;
defparam \ociram_wr_en~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(MonDReg_0),
	.datab(writedata_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.cout());
defparam \ociram_wr_data[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(address_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.cout());
defparam \ociram_addr[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_addr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[1]~1 (
	.dataa(\MonAReg[3]~q ),
	.datab(address_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.cout());
defparam \ociram_addr[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_addr[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[2]~2 (
	.dataa(\MonAReg[4]~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.cout());
defparam \ociram_addr[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_addr[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[3]~3 (
	.dataa(\MonAReg[5]~q ),
	.datab(address_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.cout());
defparam \ociram_addr[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_addr[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[4]~4 (
	.dataa(\MonAReg[6]~q ),
	.datab(address_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.cout());
defparam \ociram_addr[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_addr[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[5]~5 (
	.dataa(\MonAReg[7]~q ),
	.datab(address_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.cout());
defparam \ociram_addr[5]~5 .lut_mask = 16'hAACC;
defparam \ociram_addr[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[6]~6 (
	.dataa(\MonAReg[8]~q ),
	.datab(address_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.cout());
defparam \ociram_addr[6]~6 .lut_mask = 16'hAACC;
defparam \ociram_addr[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[7]~7 (
	.dataa(\MonAReg[9]~q ),
	.datab(address_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.cout());
defparam \ociram_addr[7]~7 .lut_mask = 16'hAACC;
defparam \ociram_addr[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.cout());
defparam \ociram_byteenable[0]~0 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(MonDReg_1),
	.datab(writedata_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.cout());
defparam \ociram_wr_data[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_wr~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_ram_wr~q ),
	.datac(jdo_35),
	.datad(\MonARegAddrInc[8]~16_combout ),
	.cin(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.cout());
defparam \jtag_ram_wr~0 .lut_mask = 16'hACFF;
defparam \jtag_ram_wr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(MonDReg_2),
	.datab(writedata_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.cout());
defparam \ociram_wr_data[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[3]~3 (
	.dataa(MonDReg_3),
	.datab(writedata_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[3]~3_combout ),
	.cout());
defparam \ociram_wr_data[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[4]~4 (
	.dataa(MonDReg_4),
	.datab(writedata_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[4]~4_combout ),
	.cout());
defparam \ociram_wr_data[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[11]~5 (
	.dataa(MonDReg_11),
	.datab(writedata_11),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[11]~5_combout ),
	.cout());
defparam \ociram_wr_data[11]~5 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[11]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[1]~1 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[1]~1_combout ),
	.cout());
defparam \ociram_byteenable[1]~1 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[13]~6 (
	.dataa(MonDReg_13),
	.datab(writedata_13),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[13]~6_combout ),
	.cout());
defparam \ociram_wr_data[13]~6 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[13]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[16]~7 (
	.dataa(MonDReg_16),
	.datab(writedata_16),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[16]~7_combout ),
	.cout());
defparam \ociram_wr_data[16]~7 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[2]~2 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[2]~2_combout ),
	.cout());
defparam \ociram_byteenable[2]~2 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[12]~8 (
	.dataa(MonDReg_12),
	.datab(writedata_12),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[12]~8_combout ),
	.cout());
defparam \ociram_wr_data[12]~8 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[12]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[5]~9 (
	.dataa(MonDReg_5),
	.datab(writedata_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[5]~9_combout ),
	.cout());
defparam \ociram_wr_data[5]~9 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[5]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[14]~10 (
	.dataa(MonDReg_14),
	.datab(writedata_14),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[14]~10_combout ),
	.cout());
defparam \ociram_wr_data[14]~10 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[14]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[15]~11 (
	.dataa(MonDReg_15),
	.datab(writedata_15),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[15]~11_combout ),
	.cout());
defparam \ociram_wr_data[15]~11 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[15]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[21]~12 (
	.dataa(MonDReg_21),
	.datab(writedata_21),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[21]~12_combout ),
	.cout());
defparam \ociram_wr_data[21]~12 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[21]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[18]~13 (
	.dataa(MonDReg_18),
	.datab(writedata_18),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[18]~13_combout ),
	.cout());
defparam \ociram_wr_data[18]~13 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[18]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[17]~14 (
	.dataa(MonDReg_17),
	.datab(writedata_17),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[17]~14_combout ),
	.cout());
defparam \ociram_wr_data[17]~14 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[17]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[31]~15 (
	.dataa(MonDReg_31),
	.datab(writedata_31),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[31]~15_combout ),
	.cout());
defparam \ociram_wr_data[31]~15 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[31]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[3]~3 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[3]~3_combout ),
	.cout());
defparam \ociram_byteenable[3]~3 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[30]~16 (
	.dataa(MonDReg_30),
	.datab(writedata_30),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[30]~16_combout ),
	.cout());
defparam \ociram_wr_data[30]~16 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[30]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[29]~17 (
	.dataa(MonDReg_29),
	.datab(writedata_29),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[29]~17_combout ),
	.cout());
defparam \ociram_wr_data[29]~17 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[29]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[28]~18 (
	.dataa(MonDReg_28),
	.datab(writedata_28),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[28]~18_combout ),
	.cout());
defparam \ociram_wr_data[28]~18 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[28]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[27]~19 (
	.dataa(MonDReg_27),
	.datab(writedata_27),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[27]~19_combout ),
	.cout());
defparam \ociram_wr_data[27]~19 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[27]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[26]~20 (
	.dataa(MonDReg_26),
	.datab(writedata_26),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[26]~20_combout ),
	.cout());
defparam \ociram_wr_data[26]~20 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[26]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[25]~21 (
	.dataa(MonDReg_25),
	.datab(writedata_25),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[25]~21_combout ),
	.cout());
defparam \ociram_wr_data[25]~21 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[25]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[10]~22 (
	.dataa(MonDReg_10),
	.datab(writedata_10),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[10]~22_combout ),
	.cout());
defparam \ociram_wr_data[10]~22 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[10]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[24]~23 (
	.dataa(MonDReg_24),
	.datab(writedata_24),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[24]~23_combout ),
	.cout());
defparam \ociram_wr_data[24]~23 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[24]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[9]~24 (
	.dataa(MonDReg_9),
	.datab(writedata_9),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[9]~24_combout ),
	.cout());
defparam \ociram_wr_data[9]~24 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[9]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[23]~25 (
	.dataa(MonDReg_23),
	.datab(writedata_23),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[23]~25_combout ),
	.cout());
defparam \ociram_wr_data[23]~25 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[8]~26 (
	.dataa(MonDReg_8),
	.datab(writedata_8),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[8]~26_combout ),
	.cout());
defparam \ociram_wr_data[8]~26 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[8]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[22]~27 (
	.dataa(MonDReg_22),
	.datab(writedata_22),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[22]~27_combout ),
	.cout());
defparam \ociram_wr_data[22]~27 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[22]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[7]~28 (
	.dataa(MonDReg_7),
	.datab(writedata_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[7]~28_combout ),
	.cout());
defparam \ociram_wr_data[7]~28 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[7]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[6]~29 (
	.dataa(MonDReg_6),
	.datab(writedata_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[6]~29_combout ),
	.cout());
defparam \ociram_wr_data[6]~29 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[6]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[20]~30 (
	.dataa(MonDReg_20),
	.datab(writedata_20),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[20]~30_combout ),
	.cout());
defparam \ociram_wr_data[20]~30 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[20]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[19]~31 (
	.dataa(MonDReg_19),
	.datab(writedata_19),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[19]~31_combout ),
	.cout());
defparam \ociram_wr_data[19]~31 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[19]~31 .sum_lutc_input = "datac";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg[0]~0_combout ),
	.asdata(jdo_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg[2]~1_combout ),
	.asdata(jdo_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg[3]~2_combout ),
	.asdata(jdo_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg[4]~3_combout ),
	.asdata(jdo_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg[29]~8_combout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(\MonDReg[28]~9_combout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[28]~24_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg[11]~5_combout ),
	.asdata(jdo_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg[12]~6_combout ),
	.asdata(jdo_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg[5]~4_combout ),
	.asdata(jdo_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg[18]~7_combout ),
	.asdata(jdo_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(\MonDReg[10]~10_combout ),
	.asdata(jdo_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~11_combout ),
	.asdata(jdo_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[28]~24_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(\MonDReg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(\MonDReg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(\MonDReg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(\MonDReg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(\MonDReg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(\MonDReg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(\MonDReg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(\MonDReg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(\MonDReg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(\MonDReg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(\MonDReg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(\MonDReg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(\MonDReg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(\MonDReg~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~12_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\MonARegAddrInc[0]~0_combout ),
	.cout(\MonARegAddrInc[0]~1 ));
defparam \MonARegAddrInc[0]~0 .lut_mask = 16'h55AA;
defparam \MonARegAddrInc[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonAReg~0 (
	.dataa(\MonARegAddrInc[0]~0_combout ),
	.datab(jdo_26),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~0_combout ),
	.cout());
defparam \MonAReg~0 .lut_mask = 16'hAACC;
defparam \MonAReg~0 .sum_lutc_input = "datac";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\MonAReg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[1]~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[0]~1 ),
	.combout(\MonARegAddrInc[1]~2_combout ),
	.cout(\MonARegAddrInc[1]~3 ));
defparam \MonARegAddrInc[1]~2 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~2 (
	.dataa(\MonARegAddrInc[1]~2_combout ),
	.datab(jdo_27),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~2_combout ),
	.cout());
defparam \MonAReg~2 .lut_mask = 16'hAACC;
defparam \MonAReg~2 .sum_lutc_input = "datac";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\MonAReg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[2]~4 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[1]~3 ),
	.combout(\MonARegAddrInc[2]~4_combout ),
	.cout(\MonARegAddrInc[2]~5 ));
defparam \MonARegAddrInc[2]~4 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~1 (
	.dataa(\MonARegAddrInc[2]~4_combout ),
	.datab(jdo_28),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~1_combout ),
	.cout());
defparam \MonAReg~1 .lut_mask = 16'hAACC;
defparam \MonAReg~1 .sum_lutc_input = "datac";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\MonAReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonAReg~3 (
	.dataa(\MonARegAddrInc[8]~16_combout ),
	.datab(jdo_17),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~3_combout ),
	.cout());
defparam \MonAReg~3 .lut_mask = 16'hAACC;
defparam \MonAReg~3 .sum_lutc_input = "datac";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\MonAReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[3]~6 (
	.dataa(\MonAReg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[2]~5 ),
	.combout(\MonARegAddrInc[3]~6_combout ),
	.cout(\MonARegAddrInc[3]~7 ));
defparam \MonARegAddrInc[3]~6 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~8 (
	.dataa(\MonARegAddrInc[3]~6_combout ),
	.datab(jdo_29),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~8_combout ),
	.cout());
defparam \MonAReg~8 .lut_mask = 16'hAACC;
defparam \MonAReg~8 .sum_lutc_input = "datac";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\MonAReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[4]~8 (
	.dataa(\MonAReg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[3]~7 ),
	.combout(\MonARegAddrInc[4]~8_combout ),
	.cout(\MonARegAddrInc[4]~9 ));
defparam \MonARegAddrInc[4]~8 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[4]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~7 (
	.dataa(\MonARegAddrInc[4]~8_combout ),
	.datab(jdo_30),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~7_combout ),
	.cout());
defparam \MonAReg~7 .lut_mask = 16'hAACC;
defparam \MonAReg~7 .sum_lutc_input = "datac";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\MonAReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[5]~10 (
	.dataa(\MonAReg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[4]~9 ),
	.combout(\MonARegAddrInc[5]~10_combout ),
	.cout(\MonARegAddrInc[5]~11 ));
defparam \MonARegAddrInc[5]~10 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~6 (
	.dataa(\MonARegAddrInc[5]~10_combout ),
	.datab(jdo_31),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~6_combout ),
	.cout());
defparam \MonAReg~6 .lut_mask = 16'hAACC;
defparam \MonAReg~6 .sum_lutc_input = "datac";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\MonAReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[6]~12 (
	.dataa(\MonAReg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[5]~11 ),
	.combout(\MonARegAddrInc[6]~12_combout ),
	.cout(\MonARegAddrInc[6]~13 ));
defparam \MonARegAddrInc[6]~12 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~5 (
	.dataa(\MonARegAddrInc[6]~12_combout ),
	.datab(jdo_32),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~5_combout ),
	.cout());
defparam \MonAReg~5 .lut_mask = 16'hAACC;
defparam \MonAReg~5 .sum_lutc_input = "datac";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\MonAReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[7]~14 (
	.dataa(\MonAReg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[6]~13 ),
	.combout(\MonARegAddrInc[7]~14_combout ),
	.cout(\MonARegAddrInc[7]~15 ));
defparam \MonARegAddrInc[7]~14 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~4 (
	.dataa(\MonARegAddrInc[7]~14_combout ),
	.datab(jdo_33),
	.datac(gnd),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\MonAReg~4_combout ),
	.cout());
defparam \MonAReg~4 .lut_mask = 16'hAACC;
defparam \MonAReg~4 .sum_lutc_input = "datac";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\MonAReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[8]~16 (
	.dataa(\MonAReg[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\MonARegAddrInc[7]~15 ),
	.combout(\MonARegAddrInc[8]~16_combout ),
	.cout());
defparam \MonARegAddrInc[8]~16 .lut_mask = 16'h5A5A;
defparam \MonARegAddrInc[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \jtag_ram_rd~0 (
	.dataa(jdo_35),
	.datab(\jtag_ram_rd~q ),
	.datac(jdo_34),
	.datad(\MonARegAddrInc[8]~16_combout ),
	.cin(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.cout());
defparam \jtag_ram_rd~0 .lut_mask = 16'hF7B3;
defparam \jtag_ram_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_rd~1 (
	.dataa(take_action_ocimem_a),
	.datab(jdo_17),
	.datac(take_action_ocimem_a1),
	.datad(\jtag_ram_rd~0_combout ),
	.cin(gnd),
	.combout(\jtag_ram_rd~1_combout ),
	.cout());
defparam \jtag_ram_rd~1 .lut_mask = 16'hFBFF;
defparam \jtag_ram_rd~1 .sum_lutc_input = "datac";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~0 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_0),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[0]~0_combout ),
	.cout());
defparam \MonDReg[0]~0 .lut_mask = 16'hAACC;
defparam \MonDReg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_rd~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_rd~q ),
	.datac(gnd),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\jtag_rd~0_combout ),
	.cout());
defparam \jtag_rd~0 .lut_mask = 16'hEEFF;
defparam \jtag_rd~0 .sum_lutc_input = "datac";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(\jtag_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~12 (
	.dataa(gnd),
	.datab(take_action_ocimem_a),
	.datac(\jtag_rd_d1~q ),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\MonDReg[0]~12_combout ),
	.cout());
defparam \MonDReg[0]~12 .lut_mask = 16'hF3C0;
defparam \MonDReg[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[2]~1 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_2),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[2]~1_combout ),
	.cout());
defparam \MonDReg[2]~1 .lut_mask = 16'hAACC;
defparam \MonDReg[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[3]~2 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_3),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[3]~2_combout ),
	.cout());
defparam \MonDReg[3]~2 .lut_mask = 16'hAACC;
defparam \MonDReg[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[4]~3 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_4),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[4]~3_combout ),
	.cout());
defparam \MonDReg[4]~3 .lut_mask = 16'hAACC;
defparam \MonDReg[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hAFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[29]~8 (
	.dataa(\Equal0~1_combout ),
	.datab(q_a_29),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[29]~8_combout ),
	.cout());
defparam \MonDReg[29]~8 .lut_mask = 16'hAACC;
defparam \MonDReg[29]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cfgrom_readdata[28]~0 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\cfgrom_readdata[28]~0_combout ),
	.cout());
defparam \cfgrom_readdata[28]~0 .lut_mask = 16'hAFFA;
defparam \cfgrom_readdata[28]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[28]~9 (
	.dataa(\cfgrom_readdata[28]~0_combout ),
	.datab(q_a_28),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[28]~9_combout ),
	.cout());
defparam \MonDReg[28]~9 .lut_mask = 16'hCC55;
defparam \MonDReg[28]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[28]~24 (
	.dataa(take_action_ocimem_b),
	.datab(\jtag_rd_d1~q ),
	.datac(gnd),
	.datad(take_action_ocimem_a),
	.cin(gnd),
	.combout(\MonDReg[28]~24_combout ),
	.cout());
defparam \MonDReg[28]~24 .lut_mask = 16'hEEFF;
defparam \MonDReg[28]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[11]~5 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_11),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[11]~5_combout ),
	.cout());
defparam \MonDReg[11]~5 .lut_mask = 16'hAACC;
defparam \MonDReg[11]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[12]~6 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_12),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[12]~6_combout ),
	.cout());
defparam \MonDReg[12]~6 .lut_mask = 16'hAACC;
defparam \MonDReg[12]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(gnd),
	.datab(\MonAReg[2]~q ),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h3FFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[5]~4 (
	.dataa(\Equal0~2_combout ),
	.datab(q_a_5),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[5]~4_combout ),
	.cout());
defparam \MonDReg[5]~4 .lut_mask = 16'hAACC;
defparam \MonDReg[5]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[2]~q ),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hAFFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[18]~7 (
	.dataa(\Equal0~3_combout ),
	.datab(q_a_18),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[18]~7_combout ),
	.cout());
defparam \MonDReg[18]~7 .lut_mask = 16'hAACC;
defparam \MonDReg[18]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[10]~10 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_10),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[10]~10_combout ),
	.cout());
defparam \MonDReg[10]~10 .lut_mask = 16'hAACC;
defparam \MonDReg[10]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cfgrom_readdata[8]~1 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\cfgrom_readdata[8]~1_combout ),
	.cout());
defparam \cfgrom_readdata[8]~1 .lut_mask = 16'hAAFF;
defparam \cfgrom_readdata[8]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[8]~11 (
	.dataa(\cfgrom_readdata[8]~1_combout ),
	.datab(q_a_8),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[8]~11_combout ),
	.cout());
defparam \MonDReg[8]~11 .lut_mask = 16'hAACC;
defparam \MonDReg[8]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~0 (
	.dataa(jdo_34),
	.datab(gnd),
	.datac(gnd),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.cout());
defparam \jtag_ram_access~0 .lut_mask = 16'hAAFF;
defparam \jtag_ram_access~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~1 (
	.dataa(jdo_17),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(\jtag_ram_access~0_combout ),
	.datad(take_action_ocimem_a),
	.cin(gnd),
	.combout(\jtag_ram_access~1_combout ),
	.cout());
defparam \jtag_ram_access~1 .lut_mask = 16'hF737;
defparam \jtag_ram_access~1 .sum_lutc_input = "datac";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cycloneive_lcell_comb \waitrequest~0 (
	.dataa(write),
	.datab(\jtag_ram_access~q ),
	.datac(address_8),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\waitrequest~0_combout ),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hEFFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(read),
	.datab(address_8),
	.datac(\jtag_ram_access~q ),
	.datad(write),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 16'hEFFF;
defparam \avalon_ociram_readdata_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~1 (
	.dataa(waitrequest1),
	.datab(\avalon_ociram_readdata_ready~0_combout ),
	.datac(write),
	.datad(\avalon_ociram_readdata_ready~q ),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~1_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~1 .lut_mask = 16'hFFFE;
defparam \avalon_ociram_readdata_ready~1 .sum_lutc_input = "datac";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cycloneive_lcell_comb \waitrequest~1 (
	.dataa(\waitrequest~0_combout ),
	.datab(read),
	.datac(\avalon_ociram_readdata_ready~q ),
	.datad(write),
	.cin(gnd),
	.combout(\waitrequest~1_combout ),
	.cout());
defparam \waitrequest~1 .lut_mask = 16'hBFFF;
defparam \waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~13 (
	.dataa(jdo_4),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_1),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~13_combout ),
	.cout());
defparam \MonDReg~13 .lut_mask = 16'hFAFC;
defparam \MonDReg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~14 (
	.dataa(jdo_19),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_16),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~14_combout ),
	.cout());
defparam \MonDReg~14 .lut_mask = 16'hFAFC;
defparam \MonDReg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~15 (
	.dataa(jdo_23),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_20),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~15_combout ),
	.cout());
defparam \MonDReg~15 .lut_mask = 16'hFAFC;
defparam \MonDReg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~16 (
	.dataa(jdo_22),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_19),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~16_combout ),
	.cout());
defparam \MonDReg~16 .lut_mask = 16'hFAFC;
defparam \MonDReg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~17 (
	.dataa(jdo_28),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_25),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~17_combout ),
	.cout());
defparam \MonDReg~17 .lut_mask = 16'hFAFC;
defparam \MonDReg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~18 (
	.dataa(jdo_30),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_27),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~18_combout ),
	.cout());
defparam \MonDReg~18 .lut_mask = 16'hFAFC;
defparam \MonDReg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~19 (
	.dataa(jdo_29),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_26),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~19_combout ),
	.cout());
defparam \MonDReg~19 .lut_mask = 16'hFAFC;
defparam \MonDReg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~20 (
	.dataa(jdo_27),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_24),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~20_combout ),
	.cout());
defparam \MonDReg~20 .lut_mask = 16'hFAFC;
defparam \MonDReg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~21 (
	.dataa(jdo_20),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_17),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~21_combout ),
	.cout());
defparam \MonDReg~21 .lut_mask = 16'hFAFC;
defparam \MonDReg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~22 (
	.dataa(jdo_34),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_31),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~22_combout ),
	.cout());
defparam \MonDReg~22 .lut_mask = 16'hFAFC;
defparam \MonDReg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~23 (
	.dataa(jdo_33),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_30),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~23_combout ),
	.cout());
defparam \MonDReg~23 .lut_mask = 16'hFAFC;
defparam \MonDReg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~25 (
	.dataa(jdo_16),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_13),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~25_combout ),
	.cout());
defparam \MonDReg~25 .lut_mask = 16'hFAFC;
defparam \MonDReg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~26 (
	.dataa(jdo_17),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_14),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~26_combout ),
	.cout());
defparam \MonDReg~26 .lut_mask = 16'hFAFC;
defparam \MonDReg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~27 (
	.dataa(jdo_18),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_15),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~27_combout ),
	.cout());
defparam \MonDReg~27 .lut_mask = 16'hFAFC;
defparam \MonDReg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~28 (
	.dataa(jdo_24),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_21),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~28_combout ),
	.cout());
defparam \MonDReg~28 .lut_mask = 16'hFAFC;
defparam \MonDReg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~29 (
	.dataa(jdo_12),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_9),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~29_combout ),
	.cout());
defparam \MonDReg~29 .lut_mask = 16'hFAFC;
defparam \MonDReg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~30 (
	.dataa(jdo_26),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_23),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~30_combout ),
	.cout());
defparam \MonDReg~30 .lut_mask = 16'hFAFC;
defparam \MonDReg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~31 (
	.dataa(jdo_25),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_22),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~31_combout ),
	.cout());
defparam \MonDReg~31 .lut_mask = 16'hFAFC;
defparam \MonDReg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~32 (
	.dataa(jdo_10),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_7),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~32_combout ),
	.cout());
defparam \MonDReg~32 .lut_mask = 16'hFAFC;
defparam \MonDReg~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~33 (
	.dataa(jdo_9),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_6),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~33_combout ),
	.cout());
defparam \MonDReg~33 .lut_mask = 16'hFAFC;
defparam \MonDReg~33 .sum_lutc_input = "datac";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_31,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_10,
	q_a_24,
	q_a_9,
	q_a_23,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	r_early_rst,
	ociram_wr_en,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_3,
	ociram_wr_data_4,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_13,
	ociram_wr_data_16,
	ociram_byteenable_2,
	ociram_wr_data_12,
	ociram_wr_data_5,
	ociram_wr_data_14,
	ociram_wr_data_15,
	ociram_wr_data_21,
	ociram_wr_data_18,
	ociram_wr_data_17,
	ociram_wr_data_31,
	ociram_byteenable_3,
	ociram_wr_data_30,
	ociram_wr_data_29,
	ociram_wr_data_28,
	ociram_wr_data_27,
	ociram_wr_data_26,
	ociram_wr_data_25,
	ociram_wr_data_10,
	ociram_wr_data_24,
	ociram_wr_data_9,
	ociram_wr_data_23,
	ociram_wr_data_8,
	ociram_wr_data_22,
	ociram_wr_data_7,
	ociram_wr_data_6,
	ociram_wr_data_20,
	ociram_wr_data_19,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_31;
output 	q_a_30;
output 	q_a_29;
output 	q_a_28;
output 	q_a_27;
output 	q_a_26;
output 	q_a_25;
output 	q_a_10;
output 	q_a_24;
output 	q_a_9;
output 	q_a_23;
output 	q_a_8;
output 	q_a_22;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_19;
input 	r_early_rst;
input 	ociram_wr_en;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_3;
input 	ociram_wr_data_4;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_13;
input 	ociram_wr_data_16;
input 	ociram_byteenable_2;
input 	ociram_wr_data_12;
input 	ociram_wr_data_5;
input 	ociram_wr_data_14;
input 	ociram_wr_data_15;
input 	ociram_wr_data_21;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	ociram_wr_data_31;
input 	ociram_byteenable_3;
input 	ociram_wr_data_30;
input 	ociram_wr_data_29;
input 	ociram_wr_data_28;
input 	ociram_wr_data_27;
input 	ociram_wr_data_26;
input 	ociram_wr_data_25;
input 	ociram_wr_data_10;
input 	ociram_wr_data_24;
input 	ociram_wr_data_9;
input 	ociram_wr_data_23;
input 	ociram_wr_data_8;
input 	ociram_wr_data_22;
input 	ociram_wr_data_7;
input 	ociram_wr_data_6;
input 	ociram_wr_data_20;
input 	ociram_wr_data_19;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(ociram_wr_en),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module final_project_soc_altsyncram_1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_4a31 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module final_project_soc_altsyncram_4a31 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_nios2_oci:the_final_project_soc_nios2_qsys_0_cpu_nios2_oci|final_project_soc_nios2_qsys_0_cpu_nios2_ocimem:the_final_project_soc_nios2_qsys_0_cpu_nios2_ocimem|final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram_module:final_project_soc_nios2_qsys_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4a31:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_register_bank_a_module (
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_31,
	q_b_30,
	q_b_29,
	D_iw_31,
	D_iw_30,
	D_iw_29,
	D_iw_28,
	D_iw_27,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_8,
	W_rf_wr_data_9,
	W_rf_wr_data_10,
	W_rf_wr_data_11,
	W_rf_wr_data_12,
	W_rf_wr_data_13,
	W_rf_wr_data_14,
	W_rf_wr_data_15,
	W_rf_wr_data_16,
	W_rf_wr_data_17,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
input 	D_iw_31;
input 	D_iw_30;
input 	D_iw_29;
input 	D_iw_28;
input 	D_iw_27;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.clock0(clk_clk));

endmodule

module final_project_soc_altsyncram_2 (
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_6mc1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module final_project_soc_altsyncram_6mc1 (
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_a_module:final_project_soc_nios2_qsys_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module final_project_soc_final_project_soc_nios2_qsys_0_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_31,
	q_b_30,
	q_b_29,
	D_iw_26,
	D_iw_25,
	D_iw_24,
	D_iw_23,
	D_iw_22,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_8,
	W_rf_wr_data_9,
	W_rf_wr_data_10,
	W_rf_wr_data_11,
	W_rf_wr_data_12,
	W_rf_wr_data_13,
	W_rf_wr_data_14,
	W_rf_wr_data_15,
	W_rf_wr_data_16,
	W_rf_wr_data_17,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_31;
output 	q_b_30;
output 	q_b_29;
input 	D_iw_26;
input 	D_iw_25;
input 	D_iw_24;
input 	D_iw_23;
input 	D_iw_22;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_3 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.clock0(clk_clk));

endmodule

module final_project_soc_altsyncram_3 (
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_6mc1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module final_project_soc_altsyncram_6mc1_1 (
	q_b,
	address_b,
	wren_a,
	data_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "final_project_soc_nios2_qsys_0:nios2_qsys_0|final_project_soc_nios2_qsys_0_cpu:cpu|final_project_soc_nios2_qsys_0_cpu_register_bank_b_module:final_project_soc_nios2_qsys_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module final_project_soc_final_project_soc_onchip_memory2_0 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_5,
	q_a_14,
	q_a_15,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_31,
	q_a_30,
	q_a_29,
	q_a_28,
	q_a_27,
	q_a_26,
	q_a_25,
	q_a_10,
	q_a_24,
	q_a_9,
	q_a_23,
	q_a_8,
	q_a_22,
	q_a_7,
	q_a_6,
	q_a_20,
	q_a_19,
	uav_write,
	saved_grant_0,
	mem_used_1,
	WideOr1,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_32,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_33,
	src_payload6,
	src_payload7,
	src_data_34,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_data_35,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_5;
output 	q_a_14;
output 	q_a_15;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_31;
output 	q_a_30;
output 	q_a_29;
output 	q_a_28;
output 	q_a_27;
output 	q_a_26;
output 	q_a_25;
output 	q_a_10;
output 	q_a_24;
output 	q_a_9;
output 	q_a_23;
output 	q_a_8;
output 	q_a_22;
output 	q_a_7;
output 	q_a_6;
output 	q_a_20;
output 	q_a_19;
input 	uav_write;
input 	saved_grant_0;
input 	mem_used_1;
input 	WideOr1;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_32;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_data_33;
input 	src_payload6;
input 	src_payload7;
input 	src_data_34;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_data_35;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


final_project_soc_altsyncram_4 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(\wren~0_combout ),
	.clocken0(r_early_rst),
	.data_a({src_payload15,src_payload16,src_payload17,src_payload18,src_payload19,src_payload20,src_payload21,src_payload23,src_payload25,src_payload27,src_payload12,src_payload30,src_payload31,src_payload13,src_payload14,src_payload7,src_payload11,src_payload10,src_payload6,
src_payload8,src_payload5,src_payload22,src_payload24,src_payload26,src_payload28,src_payload29,src_payload9,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cycloneive_lcell_comb \wren~0 (
	.dataa(mem_used_1),
	.datab(uav_write),
	.datac(saved_grant_0),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\wren~0_combout ),
	.cout());
defparam \wren~0 .lut_mask = 16'hFFFD;
defparam \wren~0 .sum_lutc_input = "datac";

endmodule

module final_project_soc_altsyncram_4 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_altsyncram_fod1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module final_project_soc_altsyncram_fod1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[1:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 2;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 3;
defparam ram_block1a0.port_a_logical_ram_depth = 4;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 2;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 3;
defparam ram_block1a1.port_a_logical_ram_depth = 4;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 2;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 3;
defparam ram_block1a2.port_a_logical_ram_depth = 4;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 2;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 3;
defparam ram_block1a3.port_a_logical_ram_depth = 4;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 2;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 3;
defparam ram_block1a4.port_a_logical_ram_depth = 4;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 2;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 3;
defparam ram_block1a11.port_a_logical_ram_depth = 4;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 2;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 3;
defparam ram_block1a13.port_a_logical_ram_depth = 4;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 2;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 3;
defparam ram_block1a16.port_a_logical_ram_depth = 4;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 2;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 3;
defparam ram_block1a12.port_a_logical_ram_depth = 4;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 2;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 3;
defparam ram_block1a5.port_a_logical_ram_depth = 4;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 2;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 3;
defparam ram_block1a14.port_a_logical_ram_depth = 4;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 2;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 3;
defparam ram_block1a15.port_a_logical_ram_depth = 4;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 2;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 3;
defparam ram_block1a21.port_a_logical_ram_depth = 4;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 2;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 3;
defparam ram_block1a18.port_a_logical_ram_depth = 4;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 2;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 3;
defparam ram_block1a17.port_a_logical_ram_depth = 4;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 2;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 3;
defparam ram_block1a31.port_a_logical_ram_depth = 4;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 2;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 3;
defparam ram_block1a30.port_a_logical_ram_depth = 4;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 2;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 3;
defparam ram_block1a29.port_a_logical_ram_depth = 4;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 2;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 3;
defparam ram_block1a28.port_a_logical_ram_depth = 4;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 2;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 3;
defparam ram_block1a27.port_a_logical_ram_depth = 4;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 2;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 3;
defparam ram_block1a26.port_a_logical_ram_depth = 4;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 2;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 3;
defparam ram_block1a25.port_a_logical_ram_depth = 4;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 2;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 3;
defparam ram_block1a10.port_a_logical_ram_depth = 4;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 2;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 3;
defparam ram_block1a24.port_a_logical_ram_depth = 4;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 2;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 3;
defparam ram_block1a9.port_a_logical_ram_depth = 4;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 2;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 3;
defparam ram_block1a23.port_a_logical_ram_depth = 4;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 2;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 3;
defparam ram_block1a8.port_a_logical_ram_depth = 4;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 2;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 3;
defparam ram_block1a22.port_a_logical_ram_depth = 4;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 2;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 3;
defparam ram_block1a7.port_a_logical_ram_depth = 4;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 2;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 3;
defparam ram_block1a6.port_a_logical_ram_depth = 4;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 2;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 3;
defparam ram_block1a20.port_a_logical_ram_depth = 4;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = 4'h0;

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "final_project_soc_onchip_memory2_0.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "final_project_soc_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_fod1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 2;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 3;
defparam ram_block1a19.port_a_logical_ram_depth = 4;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = 4'h0;

endmodule

module final_project_soc_final_project_soc_sdram (
	wire_pll7_clk_0,
	m_addr_0,
	m_addr_1,
	m_addr_2,
	m_addr_3,
	m_addr_4,
	m_addr_5,
	m_addr_6,
	m_addr_7,
	m_addr_8,
	m_addr_9,
	oe1,
	m_addr_10,
	m_addr_11,
	m_addr_12,
	m_bank_0,
	m_bank_1,
	m_cmd_1,
	m_cmd_3,
	m_dqm_0,
	m_dqm_1,
	m_dqm_2,
	m_dqm_3,
	m_cmd_2,
	m_cmd_0,
	entries_1,
	entries_0,
	altera_reset_synchronizer_int_chain_out,
	last_cycle,
	saved_grant_1,
	WideOr1,
	src_payload,
	src_data_68,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	src_data_61,
	src_data_60,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	out_data_buffer_32,
	out_data_buffer_321,
	out_data_buffer_33,
	out_data_buffer_331,
	out_data_buffer_34,
	out_data_buffer_341,
	out_data_buffer_35,
	out_data_buffer_351,
	m_data_0,
	m_data_1,
	m_data_2,
	m_data_3,
	m_data_4,
	m_data_5,
	m_data_6,
	m_data_7,
	m_data_8,
	m_data_9,
	m_data_10,
	m_data_11,
	m_data_12,
	m_data_13,
	m_data_14,
	m_data_15,
	m_data_16,
	m_data_17,
	m_data_18,
	m_data_19,
	m_data_20,
	m_data_21,
	m_data_22,
	m_data_23,
	m_data_24,
	m_data_25,
	m_data_26,
	m_data_27,
	m_data_28,
	m_data_29,
	m_data_30,
	m_data_31,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	za_valid1,
	za_data_0,
	za_data_1,
	za_data_2,
	za_data_3,
	za_data_4,
	za_data_11,
	za_data_13,
	za_data_16,
	za_data_12,
	za_data_5,
	za_data_14,
	za_data_15,
	za_data_21,
	za_data_18,
	za_data_17,
	za_data_31,
	za_data_30,
	za_data_29,
	za_data_28,
	za_data_27,
	za_data_26,
	za_data_25,
	za_data_10,
	za_data_24,
	za_data_9,
	za_data_23,
	za_data_8,
	za_data_22,
	za_data_7,
	za_data_6,
	za_data_20,
	za_data_19,
	m0_write,
	sdram_wire_dq_0,
	sdram_wire_dq_1,
	sdram_wire_dq_2,
	sdram_wire_dq_3,
	sdram_wire_dq_4,
	sdram_wire_dq_5,
	sdram_wire_dq_6,
	sdram_wire_dq_7,
	sdram_wire_dq_8,
	sdram_wire_dq_9,
	sdram_wire_dq_10,
	sdram_wire_dq_11,
	sdram_wire_dq_12,
	sdram_wire_dq_13,
	sdram_wire_dq_14,
	sdram_wire_dq_15,
	sdram_wire_dq_16,
	sdram_wire_dq_17,
	sdram_wire_dq_18,
	sdram_wire_dq_19,
	sdram_wire_dq_20,
	sdram_wire_dq_21,
	sdram_wire_dq_22,
	sdram_wire_dq_23,
	sdram_wire_dq_24,
	sdram_wire_dq_25,
	sdram_wire_dq_26,
	sdram_wire_dq_27,
	sdram_wire_dq_28,
	sdram_wire_dq_29,
	sdram_wire_dq_30,
	sdram_wire_dq_31)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_clk_0;
output 	m_addr_0;
output 	m_addr_1;
output 	m_addr_2;
output 	m_addr_3;
output 	m_addr_4;
output 	m_addr_5;
output 	m_addr_6;
output 	m_addr_7;
output 	m_addr_8;
output 	m_addr_9;
output 	oe1;
output 	m_addr_10;
output 	m_addr_11;
output 	m_addr_12;
output 	m_bank_0;
output 	m_bank_1;
output 	m_cmd_1;
output 	m_cmd_3;
output 	m_dqm_0;
output 	m_dqm_1;
output 	m_dqm_2;
output 	m_dqm_3;
output 	m_cmd_2;
output 	m_cmd_0;
output 	entries_1;
output 	entries_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	last_cycle;
input 	saved_grant_1;
input 	WideOr1;
input 	src_payload;
input 	src_data_68;
input 	src_data_48;
input 	src_data_62;
input 	src_data_49;
input 	src_data_51;
input 	src_data_50;
input 	src_data_53;
input 	src_data_52;
input 	src_data_55;
input 	src_data_54;
input 	src_data_57;
input 	src_data_56;
input 	src_data_59;
input 	src_data_58;
input 	src_data_61;
input 	src_data_60;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	out_data_buffer_32;
input 	out_data_buffer_321;
input 	out_data_buffer_33;
input 	out_data_buffer_331;
input 	out_data_buffer_34;
input 	out_data_buffer_341;
input 	out_data_buffer_35;
input 	out_data_buffer_351;
output 	m_data_0;
output 	m_data_1;
output 	m_data_2;
output 	m_data_3;
output 	m_data_4;
output 	m_data_5;
output 	m_data_6;
output 	m_data_7;
output 	m_data_8;
output 	m_data_9;
output 	m_data_10;
output 	m_data_11;
output 	m_data_12;
output 	m_data_13;
output 	m_data_14;
output 	m_data_15;
output 	m_data_16;
output 	m_data_17;
output 	m_data_18;
output 	m_data_19;
output 	m_data_20;
output 	m_data_21;
output 	m_data_22;
output 	m_data_23;
output 	m_data_24;
output 	m_data_25;
output 	m_data_26;
output 	m_data_27;
output 	m_data_28;
output 	m_data_29;
output 	m_data_30;
output 	m_data_31;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
output 	za_valid1;
output 	za_data_0;
output 	za_data_1;
output 	za_data_2;
output 	za_data_3;
output 	za_data_4;
output 	za_data_11;
output 	za_data_13;
output 	za_data_16;
output 	za_data_12;
output 	za_data_5;
output 	za_data_14;
output 	za_data_15;
output 	za_data_21;
output 	za_data_18;
output 	za_data_17;
output 	za_data_31;
output 	za_data_30;
output 	za_data_29;
output 	za_data_28;
output 	za_data_27;
output 	za_data_26;
output 	za_data_25;
output 	za_data_10;
output 	za_data_24;
output 	za_data_9;
output 	za_data_23;
output 	za_data_8;
output 	za_data_22;
output 	za_data_7;
output 	za_data_6;
output 	za_data_20;
output 	za_data_19;
input 	m0_write;
input 	sdram_wire_dq_0;
input 	sdram_wire_dq_1;
input 	sdram_wire_dq_2;
input 	sdram_wire_dq_3;
input 	sdram_wire_dq_4;
input 	sdram_wire_dq_5;
input 	sdram_wire_dq_6;
input 	sdram_wire_dq_7;
input 	sdram_wire_dq_8;
input 	sdram_wire_dq_9;
input 	sdram_wire_dq_10;
input 	sdram_wire_dq_11;
input 	sdram_wire_dq_12;
input 	sdram_wire_dq_13;
input 	sdram_wire_dq_14;
input 	sdram_wire_dq_15;
input 	sdram_wire_dq_16;
input 	sdram_wire_dq_17;
input 	sdram_wire_dq_18;
input 	sdram_wire_dq_19;
input 	sdram_wire_dq_20;
input 	sdram_wire_dq_21;
input 	sdram_wire_dq_22;
input 	sdram_wire_dq_23;
input 	sdram_wire_dq_24;
input 	sdram_wire_dq_25;
input 	sdram_wire_dq_26;
input 	sdram_wire_dq_27;
input 	sdram_wire_dq_28;
input 	sdram_wire_dq_29;
input 	sdram_wire_dq_30;
input 	sdram_wire_dq_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[46]~0_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[61]~1_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[60]~2_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[47]~3_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[49]~4_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[48]~5_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[51]~6_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[50]~7_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[53]~8_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[52]~9_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[55]~10_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[54]~11_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[57]~12_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[56]~13_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[59]~14_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[58]~15_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[36]~16_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[37]~17_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[38]~18_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[39]~19_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[40]~20_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[41]~21_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[42]~22_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[43]~23_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[44]~24_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[45]~25_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[32]~26_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[33]~27_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[34]~28_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[35]~29_combout ;
wire \comb~0_combout ;
wire \comb~1_combout ;
wire \comb~2_combout ;
wire \comb~3_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[0]~30_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[1]~31_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[2]~32_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[3]~33_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[4]~34_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[5]~35_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[6]~36_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[7]~37_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[8]~38_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[9]~39_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[10]~40_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[11]~41_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[12]~42_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[13]~43_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[14]~44_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[15]~45_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[16]~46_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[17]~47_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[18]~48_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[19]~49_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[20]~50_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[21]~51_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[22]~52_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[23]~53_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[24]~54_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[25]~55_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[26]~56_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[27]~57_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[28]~58_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[29]~59_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[30]~60_combout ;
wire \the_final_project_soc_sdram_input_efifo_module|rd_data[31]~61_combout ;
wire \Add0~0_combout ;
wire \refresh_counter~9_combout ;
wire \refresh_counter[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \refresh_counter[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \refresh_counter[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \refresh_counter~8_combout ;
wire \refresh_counter[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \refresh_counter~6_combout ;
wire \refresh_counter[4]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \refresh_counter~7_combout ;
wire \refresh_counter[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \refresh_counter~5_combout ;
wire \refresh_counter[6]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \refresh_counter[7]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \refresh_counter[8]~13_combout ;
wire \refresh_counter[8]~q ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \refresh_counter~4_combout ;
wire \refresh_counter[9]~q ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \refresh_counter~1_combout ;
wire \refresh_counter[10]~q ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \refresh_counter~3_combout ;
wire \refresh_counter[11]~q ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \refresh_counter~2_combout ;
wire \refresh_counter[12]~q ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \refresh_counter~0_combout ;
wire \refresh_counter[13]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \i_next.000~0_combout ;
wire \i_next.000~q ;
wire \Selector7~0_combout ;
wire \i_state.000~q ;
wire \Selector18~0_combout ;
wire \Selector8~0_combout ;
wire \i_state.001~q ;
wire \Selector16~0_combout ;
wire \Selector6~0_combout ;
wire \i_refs[0]~q ;
wire \Selector5~0_combout ;
wire \i_refs[1]~q ;
wire \Selector4~0_combout ;
wire \Selector4~1_combout ;
wire \i_refs[2]~q ;
wire \Selector18~1_combout ;
wire \Selector16~1_combout ;
wire \i_next.010~q ;
wire \i_count[0]~4_combout ;
wire \i_count[0]~1_combout ;
wire \i_count[0]~5_combout ;
wire \i_count[0]~q ;
wire \i_count[1]~2_combout ;
wire \i_count[1]~3_combout ;
wire \i_count[1]~q ;
wire \Selector13~0_combout ;
wire \Selector13~1_combout ;
wire \i_count[2]~q ;
wire \Selector9~0_combout ;
wire \i_state.010~q ;
wire \Selector18~2_combout ;
wire \i_next.111~q ;
wire \Selector12~0_combout ;
wire \i_state.111~q ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \i_state.011~q ;
wire \i_count[0]~0_combout ;
wire \WideOr6~0_combout ;
wire \Selector17~0_combout ;
wire \i_next.101~q ;
wire \i_state.101~0_combout ;
wire \i_state.101~q ;
wire \init_done~0_combout ;
wire \init_done~q ;
wire \Selector24~1_combout ;
wire \Selector32~0_combout ;
wire \active_rnw~q ;
wire \Selector25~5_combout ;
wire \Selector25~6_combout ;
wire \m_state.000000010~q ;
wire \active_addr[10]~q ;
wire \pending~0_combout ;
wire \active_addr[24]~q ;
wire \pending~1_combout ;
wire \active_addr[12]~q ;
wire \active_addr[13]~q ;
wire \pending~2_combout ;
wire \active_addr[14]~q ;
wire \active_addr[15]~q ;
wire \pending~3_combout ;
wire \pending~4_combout ;
wire \active_addr[16]~q ;
wire \active_addr[17]~q ;
wire \pending~5_combout ;
wire \active_addr[18]~q ;
wire \active_addr[19]~q ;
wire \pending~6_combout ;
wire \active_addr[20]~q ;
wire \active_addr[21]~q ;
wire \pending~7_combout ;
wire \active_addr[22]~q ;
wire \active_addr[23]~q ;
wire \pending~8_combout ;
wire \pending~9_combout ;
wire \m_next~19_combout ;
wire \Selector25~4_combout ;
wire \pending~10_combout ;
wire \Selector38~0_combout ;
wire \m_next~20_combout ;
wire \Selector29~0_combout ;
wire \Selector27~0_combout ;
wire \Selector35~0_combout ;
wire \Selector34~2_combout ;
wire \Selector34~3_combout ;
wire \m_next.000010000~q ;
wire \Selector27~1_combout ;
wire \Selector28~0_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \WideOr8~0_combout ;
wire \Selector27~5_combout ;
wire \Selector27~6_combout ;
wire \m_state.000010000~q ;
wire \Selector39~0_combout ;
wire \Selector39~1_combout ;
wire \Selector39~2_combout ;
wire \Selector39~3_combout ;
wire \Selector39~4_combout ;
wire \Selector39~5_combout ;
wire \m_count[0]~q ;
wire \Selector38~1_combout ;
wire \Selector38~2_combout ;
wire \Selector38~3_combout ;
wire \Selector38~4_combout ;
wire \m_count[1]~q ;
wire \Selector29~1_combout ;
wire \m_state.000100000~q ;
wire \Selector30~0_combout ;
wire \Selector30~1_combout ;
wire \m_state.001000000~q ;
wire \Selector33~0_combout ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \m_next.010000000~q ;
wire \Selector31~0_combout ;
wire \m_state.010000000~q ;
wire \Selector34~0_combout ;
wire \Selector34~1_combout ;
wire \m_next.000001000~q ;
wire \Selector27~2_combout ;
wire \m_state.000001000~q ;
wire \WideOr9~0_combout ;
wire \Selector32~1_combout ;
wire \m_state.100000000~q ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \Selector26~2_combout ;
wire \m_state.000000100~q ;
wire \Selector24~0_combout ;
wire \Selector33~1_combout ;
wire \Selector33~2_combout ;
wire \Selector33~3_combout ;
wire \Selector33~4_combout ;
wire \m_next.000000001~q ;
wire \Selector24~2_combout ;
wire \m_state.000000001~q ;
wire \Selector23~0_combout ;
wire \ack_refresh_request~q ;
wire \refresh_request~0_combout ;
wire \refresh_request~q ;
wire \active_cs_n~0_combout ;
wire \active_cs_n~1_combout ;
wire \active_cs_n~q ;
wire \pending~combout ;
wire \active_rnw~2_combout ;
wire \active_rnw~4_combout ;
wire \active_rnw~3_combout ;
wire \active_addr[11]~q ;
wire \Selector41~0_combout ;
wire \Selector41~1_combout ;
wire \f_pop~q ;
wire \m_addr[3]~0_combout ;
wire \active_addr[0]~q ;
wire \i_addr[12]~q ;
wire \Selector116~0_combout ;
wire \Selector116~1_combout ;
wire \m_addr[3]~1_combout ;
wire \m_addr[3]~2_combout ;
wire \active_addr[1]~q ;
wire \Selector115~0_combout ;
wire \Selector115~1_combout ;
wire \active_addr[2]~q ;
wire \Selector114~0_combout ;
wire \Selector114~1_combout ;
wire \active_addr[3]~q ;
wire \Selector113~0_combout ;
wire \Selector113~1_combout ;
wire \active_addr[4]~q ;
wire \Selector112~0_combout ;
wire \Selector112~1_combout ;
wire \active_addr[5]~q ;
wire \f_select~combout ;
wire \Selector111~0_combout ;
wire \Selector111~1_combout ;
wire \active_addr[6]~q ;
wire \Selector110~0_combout ;
wire \Selector110~1_combout ;
wire \active_addr[7]~q ;
wire \Selector109~0_combout ;
wire \Selector109~1_combout ;
wire \active_addr[8]~q ;
wire \Selector108~0_combout ;
wire \Selector108~1_combout ;
wire \active_addr[9]~q ;
wire \Selector107~0_combout ;
wire \Selector107~1_combout ;
wire \always5~0_combout ;
wire \Selector106~2_combout ;
wire \Selector106~3_combout ;
wire \Selector105~2_combout ;
wire \Selector105~3_combout ;
wire \Selector104~2_combout ;
wire \Selector104~3_combout ;
wire \Selector118~0_combout ;
wire \WideOr16~0_combout ;
wire \Selector117~0_combout ;
wire \Selector2~0_combout ;
wire \i_cmd[1]~q ;
wire \Selector21~0_combout ;
wire \Selector21~1_combout ;
wire \Selector0~0_combout ;
wire \i_cmd[3]~q ;
wire \Selector19~0_combout ;
wire \Selector19~1_combout ;
wire \Selector19~2_combout ;
wire \Selector19~3_combout ;
wire \active_dqm[0]~q ;
wire \Selector154~0_combout ;
wire \active_dqm[1]~q ;
wire \Selector153~0_combout ;
wire \active_dqm[2]~q ;
wire \Selector152~0_combout ;
wire \active_dqm[3]~q ;
wire \Selector151~0_combout ;
wire \Selector1~0_combout ;
wire \i_cmd[2]~q ;
wire \Selector20~0_combout ;
wire \Selector3~0_combout ;
wire \i_cmd[0]~q ;
wire \Selector22~0_combout ;
wire \Selector22~1_combout ;
wire \active_data[0]~q ;
wire \Selector150~0_combout ;
wire \m_data[3]~0_combout ;
wire \Selector150~1_combout ;
wire \active_data[1]~q ;
wire \Selector149~0_combout ;
wire \Selector149~1_combout ;
wire \active_data[2]~q ;
wire \Selector148~0_combout ;
wire \Selector148~1_combout ;
wire \active_data[3]~q ;
wire \Selector147~0_combout ;
wire \Selector147~1_combout ;
wire \active_data[4]~q ;
wire \Selector146~0_combout ;
wire \Selector146~1_combout ;
wire \active_data[5]~q ;
wire \Selector145~0_combout ;
wire \Selector145~1_combout ;
wire \active_data[6]~q ;
wire \Selector144~0_combout ;
wire \Selector144~1_combout ;
wire \active_data[7]~q ;
wire \Selector143~0_combout ;
wire \Selector143~1_combout ;
wire \active_data[8]~q ;
wire \Selector142~0_combout ;
wire \Selector142~1_combout ;
wire \active_data[9]~q ;
wire \Selector141~0_combout ;
wire \Selector141~1_combout ;
wire \active_data[10]~q ;
wire \Selector140~0_combout ;
wire \Selector140~1_combout ;
wire \active_data[11]~q ;
wire \Selector139~0_combout ;
wire \Selector139~1_combout ;
wire \active_data[12]~q ;
wire \Selector138~0_combout ;
wire \Selector138~1_combout ;
wire \active_data[13]~q ;
wire \Selector137~0_combout ;
wire \Selector137~1_combout ;
wire \active_data[14]~q ;
wire \Selector136~0_combout ;
wire \Selector136~1_combout ;
wire \active_data[15]~q ;
wire \Selector135~0_combout ;
wire \Selector135~1_combout ;
wire \active_data[16]~q ;
wire \Selector134~0_combout ;
wire \Selector134~1_combout ;
wire \active_data[17]~q ;
wire \Selector133~0_combout ;
wire \Selector133~1_combout ;
wire \active_data[18]~q ;
wire \Selector132~0_combout ;
wire \Selector132~1_combout ;
wire \active_data[19]~q ;
wire \Selector131~0_combout ;
wire \Selector131~1_combout ;
wire \active_data[20]~q ;
wire \Selector130~0_combout ;
wire \Selector130~1_combout ;
wire \active_data[21]~q ;
wire \Selector129~0_combout ;
wire \Selector129~1_combout ;
wire \active_data[22]~q ;
wire \Selector128~0_combout ;
wire \Selector128~1_combout ;
wire \active_data[23]~q ;
wire \Selector127~0_combout ;
wire \Selector127~1_combout ;
wire \active_data[24]~q ;
wire \Selector126~0_combout ;
wire \Selector126~1_combout ;
wire \active_data[25]~q ;
wire \Selector125~0_combout ;
wire \Selector125~1_combout ;
wire \active_data[26]~q ;
wire \Selector124~0_combout ;
wire \Selector124~1_combout ;
wire \active_data[27]~q ;
wire \Selector123~0_combout ;
wire \Selector123~1_combout ;
wire \active_data[28]~q ;
wire \Selector122~0_combout ;
wire \Selector122~1_combout ;
wire \active_data[29]~q ;
wire \Selector121~0_combout ;
wire \Selector121~1_combout ;
wire \active_data[30]~q ;
wire \Selector120~0_combout ;
wire \Selector120~1_combout ;
wire \active_data[31]~q ;
wire \Selector119~0_combout ;
wire \Selector119~1_combout ;
wire \Equal4~0_combout ;
wire \rd_valid[0]~q ;
wire \rd_valid[1]~q ;
wire \rd_valid[2]~q ;


final_project_soc_final_project_soc_sdram_input_efifo_module the_final_project_soc_sdram_input_efifo_module(
	.clk(wire_pll7_clk_0),
	.f_pop(\f_pop~q ),
	.entries_1(entries_1),
	.entries_0(entries_0),
	.Equal1(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.rd_data_46(\the_final_project_soc_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.rd_data_61(\the_final_project_soc_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.rd_data_60(\the_final_project_soc_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.rd_data_47(\the_final_project_soc_sdram_input_efifo_module|rd_data[47]~3_combout ),
	.rd_data_49(\the_final_project_soc_sdram_input_efifo_module|rd_data[49]~4_combout ),
	.rd_data_48(\the_final_project_soc_sdram_input_efifo_module|rd_data[48]~5_combout ),
	.rd_data_51(\the_final_project_soc_sdram_input_efifo_module|rd_data[51]~6_combout ),
	.rd_data_50(\the_final_project_soc_sdram_input_efifo_module|rd_data[50]~7_combout ),
	.rd_data_53(\the_final_project_soc_sdram_input_efifo_module|rd_data[53]~8_combout ),
	.rd_data_52(\the_final_project_soc_sdram_input_efifo_module|rd_data[52]~9_combout ),
	.rd_data_55(\the_final_project_soc_sdram_input_efifo_module|rd_data[55]~10_combout ),
	.rd_data_54(\the_final_project_soc_sdram_input_efifo_module|rd_data[54]~11_combout ),
	.rd_data_57(\the_final_project_soc_sdram_input_efifo_module|rd_data[57]~12_combout ),
	.rd_data_56(\the_final_project_soc_sdram_input_efifo_module|rd_data[56]~13_combout ),
	.rd_data_59(\the_final_project_soc_sdram_input_efifo_module|rd_data[59]~14_combout ),
	.rd_data_58(\the_final_project_soc_sdram_input_efifo_module|rd_data[58]~15_combout ),
	.pending(\pending~combout ),
	.rd_data_36(\the_final_project_soc_sdram_input_efifo_module|rd_data[36]~16_combout ),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.rd_data_37(\the_final_project_soc_sdram_input_efifo_module|rd_data[37]~17_combout ),
	.rd_data_38(\the_final_project_soc_sdram_input_efifo_module|rd_data[38]~18_combout ),
	.rd_data_39(\the_final_project_soc_sdram_input_efifo_module|rd_data[39]~19_combout ),
	.rd_data_40(\the_final_project_soc_sdram_input_efifo_module|rd_data[40]~20_combout ),
	.rd_data_41(\the_final_project_soc_sdram_input_efifo_module|rd_data[41]~21_combout ),
	.f_select(\f_select~combout ),
	.rd_data_42(\the_final_project_soc_sdram_input_efifo_module|rd_data[42]~22_combout ),
	.rd_data_43(\the_final_project_soc_sdram_input_efifo_module|rd_data[43]~23_combout ),
	.rd_data_44(\the_final_project_soc_sdram_input_efifo_module|rd_data[44]~24_combout ),
	.rd_data_45(\the_final_project_soc_sdram_input_efifo_module|rd_data[45]~25_combout ),
	.rd_data_32(\the_final_project_soc_sdram_input_efifo_module|rd_data[32]~26_combout ),
	.rd_data_33(\the_final_project_soc_sdram_input_efifo_module|rd_data[33]~27_combout ),
	.rd_data_34(\the_final_project_soc_sdram_input_efifo_module|rd_data[34]~28_combout ),
	.rd_data_35(\the_final_project_soc_sdram_input_efifo_module|rd_data[35]~29_combout ),
	.last_cycle(last_cycle),
	.WideOr1(WideOr1),
	.src_payload(src_payload),
	.src_data_68(src_data_68),
	.src_data_48(src_data_48),
	.src_data_62(src_data_62),
	.src_data_49(src_data_49),
	.src_data_51(src_data_51),
	.src_data_50(src_data_50),
	.src_data_53(src_data_53),
	.src_data_52(src_data_52),
	.src_data_55(src_data_55),
	.src_data_54(src_data_54),
	.src_data_57(src_data_57),
	.src_data_56(src_data_56),
	.src_data_59(src_data_59),
	.src_data_58(src_data_58),
	.src_data_61(src_data_61),
	.src_data_60(src_data_60),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_46),
	.src_data_47(src_data_47),
	.comb(\comb~0_combout ),
	.comb1(\comb~1_combout ),
	.comb2(\comb~2_combout ),
	.comb3(\comb~3_combout ),
	.rd_data_0(\the_final_project_soc_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.rd_data_1(\the_final_project_soc_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.rd_data_2(\the_final_project_soc_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.rd_data_3(\the_final_project_soc_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.rd_data_4(\the_final_project_soc_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.rd_data_5(\the_final_project_soc_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.rd_data_6(\the_final_project_soc_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.rd_data_7(\the_final_project_soc_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.rd_data_8(\the_final_project_soc_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.rd_data_9(\the_final_project_soc_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.rd_data_10(\the_final_project_soc_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.rd_data_11(\the_final_project_soc_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.rd_data_12(\the_final_project_soc_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.rd_data_13(\the_final_project_soc_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.rd_data_14(\the_final_project_soc_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.rd_data_15(\the_final_project_soc_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.rd_data_16(\the_final_project_soc_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.rd_data_17(\the_final_project_soc_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.rd_data_18(\the_final_project_soc_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.rd_data_19(\the_final_project_soc_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.rd_data_20(\the_final_project_soc_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.rd_data_21(\the_final_project_soc_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.rd_data_22(\the_final_project_soc_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.rd_data_23(\the_final_project_soc_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.rd_data_24(\the_final_project_soc_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.rd_data_25(\the_final_project_soc_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.rd_data_26(\the_final_project_soc_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.rd_data_27(\the_final_project_soc_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.rd_data_28(\the_final_project_soc_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.rd_data_29(\the_final_project_soc_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.rd_data_30(\the_final_project_soc_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.rd_data_31(\the_final_project_soc_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.m0_write(m0_write));

cycloneive_lcell_comb \comb~0 (
	.dataa(out_data_buffer_32),
	.datab(saved_grant_1),
	.datac(out_data_buffer_321),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'h7FFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~1 (
	.dataa(out_data_buffer_33),
	.datab(saved_grant_1),
	.datac(out_data_buffer_331),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'h7FFF;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~2 (
	.dataa(out_data_buffer_34),
	.datab(saved_grant_1),
	.datac(out_data_buffer_341),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
defparam \comb~2 .lut_mask = 16'h7FFF;
defparam \comb~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~3 (
	.dataa(out_data_buffer_35),
	.datab(saved_grant_1),
	.datac(out_data_buffer_351),
	.datad(m0_write),
	.cin(gnd),
	.combout(\comb~3_combout ),
	.cout());
defparam \comb~3 .lut_mask = 16'h7FFF;
defparam \comb~3 .sum_lutc_input = "datac";

dffeas \m_addr[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector116~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_0),
	.prn(vcc));
defparam \m_addr[0] .is_wysiwyg = "true";
defparam \m_addr[0] .power_up = "low";

dffeas \m_addr[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector115~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_1),
	.prn(vcc));
defparam \m_addr[1] .is_wysiwyg = "true";
defparam \m_addr[1] .power_up = "low";

dffeas \m_addr[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector114~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_2),
	.prn(vcc));
defparam \m_addr[2] .is_wysiwyg = "true";
defparam \m_addr[2] .power_up = "low";

dffeas \m_addr[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector113~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_3),
	.prn(vcc));
defparam \m_addr[3] .is_wysiwyg = "true";
defparam \m_addr[3] .power_up = "low";

dffeas \m_addr[4] (
	.clk(wire_pll7_clk_0),
	.d(\Selector112~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_4),
	.prn(vcc));
defparam \m_addr[4] .is_wysiwyg = "true";
defparam \m_addr[4] .power_up = "low";

dffeas \m_addr[5] (
	.clk(wire_pll7_clk_0),
	.d(\Selector111~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_5),
	.prn(vcc));
defparam \m_addr[5] .is_wysiwyg = "true";
defparam \m_addr[5] .power_up = "low";

dffeas \m_addr[6] (
	.clk(wire_pll7_clk_0),
	.d(\Selector110~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_6),
	.prn(vcc));
defparam \m_addr[6] .is_wysiwyg = "true";
defparam \m_addr[6] .power_up = "low";

dffeas \m_addr[7] (
	.clk(wire_pll7_clk_0),
	.d(\Selector109~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_7),
	.prn(vcc));
defparam \m_addr[7] .is_wysiwyg = "true";
defparam \m_addr[7] .power_up = "low";

dffeas \m_addr[8] (
	.clk(wire_pll7_clk_0),
	.d(\Selector108~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_8),
	.prn(vcc));
defparam \m_addr[8] .is_wysiwyg = "true";
defparam \m_addr[8] .power_up = "low";

dffeas \m_addr[9] (
	.clk(wire_pll7_clk_0),
	.d(\Selector107~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\m_state.001000000~q ),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_9),
	.prn(vcc));
defparam \m_addr[9] .is_wysiwyg = "true";
defparam \m_addr[9] .power_up = "low";

dffeas oe(
	.clk(wire_pll7_clk_0),
	.d(\always5~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(!\m_state.000010000~q ),
	.sload(gnd),
	.ena(vcc),
	.q(oe1),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

dffeas \m_addr[10] (
	.clk(wire_pll7_clk_0),
	.d(\Selector106~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_10),
	.prn(vcc));
defparam \m_addr[10] .is_wysiwyg = "true";
defparam \m_addr[10] .power_up = "low";

dffeas \m_addr[11] (
	.clk(wire_pll7_clk_0),
	.d(\Selector105~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_11),
	.prn(vcc));
defparam \m_addr[11] .is_wysiwyg = "true";
defparam \m_addr[11] .power_up = "low";

dffeas \m_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\Selector104~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\m_addr[3]~2_combout ),
	.q(m_addr_12),
	.prn(vcc));
defparam \m_addr[12] .is_wysiwyg = "true";
defparam \m_addr[12] .power_up = "low";

dffeas \m_bank[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector118~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_0),
	.prn(vcc));
defparam \m_bank[0] .is_wysiwyg = "true";
defparam \m_bank[0] .power_up = "low";

dffeas \m_bank[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector117~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_bank_1),
	.prn(vcc));
defparam \m_bank[1] .is_wysiwyg = "true";
defparam \m_bank[1] .power_up = "low";

dffeas \m_cmd[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector21~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_1),
	.prn(vcc));
defparam \m_cmd[1] .is_wysiwyg = "true";
defparam \m_cmd[1] .power_up = "low";

dffeas \m_cmd[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector19~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_3),
	.prn(vcc));
defparam \m_cmd[3] .is_wysiwyg = "true";
defparam \m_cmd[3] .power_up = "low";

dffeas \m_dqm[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector154~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_0),
	.prn(vcc));
defparam \m_dqm[0] .is_wysiwyg = "true";
defparam \m_dqm[0] .power_up = "low";

dffeas \m_dqm[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector153~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_1),
	.prn(vcc));
defparam \m_dqm[1] .is_wysiwyg = "true";
defparam \m_dqm[1] .power_up = "low";

dffeas \m_dqm[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector152~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_2),
	.prn(vcc));
defparam \m_dqm[2] .is_wysiwyg = "true";
defparam \m_dqm[2] .power_up = "low";

dffeas \m_dqm[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector151~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WideOr16~0_combout ),
	.q(m_dqm_3),
	.prn(vcc));
defparam \m_dqm[3] .is_wysiwyg = "true";
defparam \m_dqm[3] .power_up = "low";

dffeas \m_cmd[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_2),
	.prn(vcc));
defparam \m_cmd[2] .is_wysiwyg = "true";
defparam \m_cmd[2] .power_up = "low";

dffeas \m_cmd[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector22~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_cmd_0),
	.prn(vcc));
defparam \m_cmd[0] .is_wysiwyg = "true";
defparam \m_cmd[0] .power_up = "low";

dffeas \m_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector150~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_0),
	.prn(vcc));
defparam \m_data[0] .is_wysiwyg = "true";
defparam \m_data[0] .power_up = "low";

dffeas \m_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector149~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_1),
	.prn(vcc));
defparam \m_data[1] .is_wysiwyg = "true";
defparam \m_data[1] .power_up = "low";

dffeas \m_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector148~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_2),
	.prn(vcc));
defparam \m_data[2] .is_wysiwyg = "true";
defparam \m_data[2] .power_up = "low";

dffeas \m_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector147~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_3),
	.prn(vcc));
defparam \m_data[3] .is_wysiwyg = "true";
defparam \m_data[3] .power_up = "low";

dffeas \m_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\Selector146~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_4),
	.prn(vcc));
defparam \m_data[4] .is_wysiwyg = "true";
defparam \m_data[4] .power_up = "low";

dffeas \m_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\Selector145~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_5),
	.prn(vcc));
defparam \m_data[5] .is_wysiwyg = "true";
defparam \m_data[5] .power_up = "low";

dffeas \m_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\Selector144~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_6),
	.prn(vcc));
defparam \m_data[6] .is_wysiwyg = "true";
defparam \m_data[6] .power_up = "low";

dffeas \m_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\Selector143~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_7),
	.prn(vcc));
defparam \m_data[7] .is_wysiwyg = "true";
defparam \m_data[7] .power_up = "low";

dffeas \m_data[8] (
	.clk(wire_pll7_clk_0),
	.d(\Selector142~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_8),
	.prn(vcc));
defparam \m_data[8] .is_wysiwyg = "true";
defparam \m_data[8] .power_up = "low";

dffeas \m_data[9] (
	.clk(wire_pll7_clk_0),
	.d(\Selector141~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_9),
	.prn(vcc));
defparam \m_data[9] .is_wysiwyg = "true";
defparam \m_data[9] .power_up = "low";

dffeas \m_data[10] (
	.clk(wire_pll7_clk_0),
	.d(\Selector140~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_10),
	.prn(vcc));
defparam \m_data[10] .is_wysiwyg = "true";
defparam \m_data[10] .power_up = "low";

dffeas \m_data[11] (
	.clk(wire_pll7_clk_0),
	.d(\Selector139~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_11),
	.prn(vcc));
defparam \m_data[11] .is_wysiwyg = "true";
defparam \m_data[11] .power_up = "low";

dffeas \m_data[12] (
	.clk(wire_pll7_clk_0),
	.d(\Selector138~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_12),
	.prn(vcc));
defparam \m_data[12] .is_wysiwyg = "true";
defparam \m_data[12] .power_up = "low";

dffeas \m_data[13] (
	.clk(wire_pll7_clk_0),
	.d(\Selector137~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_13),
	.prn(vcc));
defparam \m_data[13] .is_wysiwyg = "true";
defparam \m_data[13] .power_up = "low";

dffeas \m_data[14] (
	.clk(wire_pll7_clk_0),
	.d(\Selector136~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_14),
	.prn(vcc));
defparam \m_data[14] .is_wysiwyg = "true";
defparam \m_data[14] .power_up = "low";

dffeas \m_data[15] (
	.clk(wire_pll7_clk_0),
	.d(\Selector135~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_15),
	.prn(vcc));
defparam \m_data[15] .is_wysiwyg = "true";
defparam \m_data[15] .power_up = "low";

dffeas \m_data[16] (
	.clk(wire_pll7_clk_0),
	.d(\Selector134~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_16),
	.prn(vcc));
defparam \m_data[16] .is_wysiwyg = "true";
defparam \m_data[16] .power_up = "low";

dffeas \m_data[17] (
	.clk(wire_pll7_clk_0),
	.d(\Selector133~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_17),
	.prn(vcc));
defparam \m_data[17] .is_wysiwyg = "true";
defparam \m_data[17] .power_up = "low";

dffeas \m_data[18] (
	.clk(wire_pll7_clk_0),
	.d(\Selector132~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_18),
	.prn(vcc));
defparam \m_data[18] .is_wysiwyg = "true";
defparam \m_data[18] .power_up = "low";

dffeas \m_data[19] (
	.clk(wire_pll7_clk_0),
	.d(\Selector131~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_19),
	.prn(vcc));
defparam \m_data[19] .is_wysiwyg = "true";
defparam \m_data[19] .power_up = "low";

dffeas \m_data[20] (
	.clk(wire_pll7_clk_0),
	.d(\Selector130~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_20),
	.prn(vcc));
defparam \m_data[20] .is_wysiwyg = "true";
defparam \m_data[20] .power_up = "low";

dffeas \m_data[21] (
	.clk(wire_pll7_clk_0),
	.d(\Selector129~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_21),
	.prn(vcc));
defparam \m_data[21] .is_wysiwyg = "true";
defparam \m_data[21] .power_up = "low";

dffeas \m_data[22] (
	.clk(wire_pll7_clk_0),
	.d(\Selector128~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_22),
	.prn(vcc));
defparam \m_data[22] .is_wysiwyg = "true";
defparam \m_data[22] .power_up = "low";

dffeas \m_data[23] (
	.clk(wire_pll7_clk_0),
	.d(\Selector127~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_23),
	.prn(vcc));
defparam \m_data[23] .is_wysiwyg = "true";
defparam \m_data[23] .power_up = "low";

dffeas \m_data[24] (
	.clk(wire_pll7_clk_0),
	.d(\Selector126~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_24),
	.prn(vcc));
defparam \m_data[24] .is_wysiwyg = "true";
defparam \m_data[24] .power_up = "low";

dffeas \m_data[25] (
	.clk(wire_pll7_clk_0),
	.d(\Selector125~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_25),
	.prn(vcc));
defparam \m_data[25] .is_wysiwyg = "true";
defparam \m_data[25] .power_up = "low";

dffeas \m_data[26] (
	.clk(wire_pll7_clk_0),
	.d(\Selector124~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_26),
	.prn(vcc));
defparam \m_data[26] .is_wysiwyg = "true";
defparam \m_data[26] .power_up = "low";

dffeas \m_data[27] (
	.clk(wire_pll7_clk_0),
	.d(\Selector123~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_27),
	.prn(vcc));
defparam \m_data[27] .is_wysiwyg = "true";
defparam \m_data[27] .power_up = "low";

dffeas \m_data[28] (
	.clk(wire_pll7_clk_0),
	.d(\Selector122~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_28),
	.prn(vcc));
defparam \m_data[28] .is_wysiwyg = "true";
defparam \m_data[28] .power_up = "low";

dffeas \m_data[29] (
	.clk(wire_pll7_clk_0),
	.d(\Selector121~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_29),
	.prn(vcc));
defparam \m_data[29] .is_wysiwyg = "true";
defparam \m_data[29] .power_up = "low";

dffeas \m_data[30] (
	.clk(wire_pll7_clk_0),
	.d(\Selector120~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_30),
	.prn(vcc));
defparam \m_data[30] .is_wysiwyg = "true";
defparam \m_data[30] .power_up = "low";

dffeas \m_data[31] (
	.clk(wire_pll7_clk_0),
	.d(\Selector119~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(m_data_31),
	.prn(vcc));
defparam \m_data[31] .is_wysiwyg = "true";
defparam \m_data[31] .power_up = "low";

dffeas za_valid(
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[2]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_valid1),
	.prn(vcc));
defparam za_valid.is_wysiwyg = "true";
defparam za_valid.power_up = "low";

dffeas \za_data[0] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_0),
	.prn(vcc));
defparam \za_data[0] .is_wysiwyg = "true";
defparam \za_data[0] .power_up = "low";

dffeas \za_data[1] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_1),
	.prn(vcc));
defparam \za_data[1] .is_wysiwyg = "true";
defparam \za_data[1] .power_up = "low";

dffeas \za_data[2] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_2),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_2),
	.prn(vcc));
defparam \za_data[2] .is_wysiwyg = "true";
defparam \za_data[2] .power_up = "low";

dffeas \za_data[3] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_3),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_3),
	.prn(vcc));
defparam \za_data[3] .is_wysiwyg = "true";
defparam \za_data[3] .power_up = "low";

dffeas \za_data[4] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_4),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_4),
	.prn(vcc));
defparam \za_data[4] .is_wysiwyg = "true";
defparam \za_data[4] .power_up = "low";

dffeas \za_data[11] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_11),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_11),
	.prn(vcc));
defparam \za_data[11] .is_wysiwyg = "true";
defparam \za_data[11] .power_up = "low";

dffeas \za_data[13] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_13),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_13),
	.prn(vcc));
defparam \za_data[13] .is_wysiwyg = "true";
defparam \za_data[13] .power_up = "low";

dffeas \za_data[16] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_16),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_16),
	.prn(vcc));
defparam \za_data[16] .is_wysiwyg = "true";
defparam \za_data[16] .power_up = "low";

dffeas \za_data[12] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_12),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_12),
	.prn(vcc));
defparam \za_data[12] .is_wysiwyg = "true";
defparam \za_data[12] .power_up = "low";

dffeas \za_data[5] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_5),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_5),
	.prn(vcc));
defparam \za_data[5] .is_wysiwyg = "true";
defparam \za_data[5] .power_up = "low";

dffeas \za_data[14] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_14),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_14),
	.prn(vcc));
defparam \za_data[14] .is_wysiwyg = "true";
defparam \za_data[14] .power_up = "low";

dffeas \za_data[15] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_15),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_15),
	.prn(vcc));
defparam \za_data[15] .is_wysiwyg = "true";
defparam \za_data[15] .power_up = "low";

dffeas \za_data[21] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_21),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_21),
	.prn(vcc));
defparam \za_data[21] .is_wysiwyg = "true";
defparam \za_data[21] .power_up = "low";

dffeas \za_data[18] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_18),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_18),
	.prn(vcc));
defparam \za_data[18] .is_wysiwyg = "true";
defparam \za_data[18] .power_up = "low";

dffeas \za_data[17] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_17),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_17),
	.prn(vcc));
defparam \za_data[17] .is_wysiwyg = "true";
defparam \za_data[17] .power_up = "low";

dffeas \za_data[31] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_31),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_31),
	.prn(vcc));
defparam \za_data[31] .is_wysiwyg = "true";
defparam \za_data[31] .power_up = "low";

dffeas \za_data[30] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_30),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_30),
	.prn(vcc));
defparam \za_data[30] .is_wysiwyg = "true";
defparam \za_data[30] .power_up = "low";

dffeas \za_data[29] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_29),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_29),
	.prn(vcc));
defparam \za_data[29] .is_wysiwyg = "true";
defparam \za_data[29] .power_up = "low";

dffeas \za_data[28] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_28),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_28),
	.prn(vcc));
defparam \za_data[28] .is_wysiwyg = "true";
defparam \za_data[28] .power_up = "low";

dffeas \za_data[27] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_27),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_27),
	.prn(vcc));
defparam \za_data[27] .is_wysiwyg = "true";
defparam \za_data[27] .power_up = "low";

dffeas \za_data[26] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_26),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_26),
	.prn(vcc));
defparam \za_data[26] .is_wysiwyg = "true";
defparam \za_data[26] .power_up = "low";

dffeas \za_data[25] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_25),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_25),
	.prn(vcc));
defparam \za_data[25] .is_wysiwyg = "true";
defparam \za_data[25] .power_up = "low";

dffeas \za_data[10] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_10),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_10),
	.prn(vcc));
defparam \za_data[10] .is_wysiwyg = "true";
defparam \za_data[10] .power_up = "low";

dffeas \za_data[24] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_24),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_24),
	.prn(vcc));
defparam \za_data[24] .is_wysiwyg = "true";
defparam \za_data[24] .power_up = "low";

dffeas \za_data[9] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_9),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_9),
	.prn(vcc));
defparam \za_data[9] .is_wysiwyg = "true";
defparam \za_data[9] .power_up = "low";

dffeas \za_data[23] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_23),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_23),
	.prn(vcc));
defparam \za_data[23] .is_wysiwyg = "true";
defparam \za_data[23] .power_up = "low";

dffeas \za_data[8] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_8),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_8),
	.prn(vcc));
defparam \za_data[8] .is_wysiwyg = "true";
defparam \za_data[8] .power_up = "low";

dffeas \za_data[22] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_22),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_22),
	.prn(vcc));
defparam \za_data[22] .is_wysiwyg = "true";
defparam \za_data[22] .power_up = "low";

dffeas \za_data[7] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_7),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_7),
	.prn(vcc));
defparam \za_data[7] .is_wysiwyg = "true";
defparam \za_data[7] .power_up = "low";

dffeas \za_data[6] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_6),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_6),
	.prn(vcc));
defparam \za_data[6] .is_wysiwyg = "true";
defparam \za_data[6] .power_up = "low";

dffeas \za_data[20] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_20),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_20),
	.prn(vcc));
defparam \za_data[20] .is_wysiwyg = "true";
defparam \za_data[20] .power_up = "low";

dffeas \za_data[19] (
	.clk(wire_pll7_clk_0),
	.d(sdram_wire_dq_19),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(za_data_19),
	.prn(vcc));
defparam \za_data[19] .is_wysiwyg = "true";
defparam \za_data[19] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\refresh_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \refresh_counter~9 (
	.dataa(\Add0~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~9_combout ),
	.cout());
defparam \refresh_counter~9 .lut_mask = 16'hAAFF;
defparam \refresh_counter~9 .sum_lutc_input = "datac";

dffeas \refresh_counter[0] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[0]~q ),
	.prn(vcc));
defparam \refresh_counter[0] .is_wysiwyg = "true";
defparam \refresh_counter[0] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\refresh_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

dffeas \refresh_counter[1] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[1]~q ),
	.prn(vcc));
defparam \refresh_counter[1] .is_wysiwyg = "true";
defparam \refresh_counter[1] .power_up = "low";

cycloneive_lcell_comb \Add0~4 (
	.dataa(\refresh_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

dffeas \refresh_counter[2] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[2]~q ),
	.prn(vcc));
defparam \refresh_counter[2] .is_wysiwyg = "true";
defparam \refresh_counter[2] .power_up = "low";

cycloneive_lcell_comb \Add0~6 (
	.dataa(\refresh_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~8 (
	.dataa(\Add0~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~8_combout ),
	.cout());
defparam \refresh_counter~8 .lut_mask = 16'hAAFF;
defparam \refresh_counter~8 .sum_lutc_input = "datac";

dffeas \refresh_counter[3] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[3]~q ),
	.prn(vcc));
defparam \refresh_counter[3] .is_wysiwyg = "true";
defparam \refresh_counter[3] .power_up = "low";

cycloneive_lcell_comb \Add0~8 (
	.dataa(\refresh_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~6 (
	.dataa(\Add0~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~6_combout ),
	.cout());
defparam \refresh_counter~6 .lut_mask = 16'hFF55;
defparam \refresh_counter~6 .sum_lutc_input = "datac";

dffeas \refresh_counter[4] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[4]~q ),
	.prn(vcc));
defparam \refresh_counter[4] .is_wysiwyg = "true";
defparam \refresh_counter[4] .power_up = "low";

cycloneive_lcell_comb \Add0~10 (
	.dataa(\refresh_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~7 (
	.dataa(\Add0~10_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~7_combout ),
	.cout());
defparam \refresh_counter~7 .lut_mask = 16'hAAFF;
defparam \refresh_counter~7 .sum_lutc_input = "datac";

dffeas \refresh_counter[5] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[5]~q ),
	.prn(vcc));
defparam \refresh_counter[5] .is_wysiwyg = "true";
defparam \refresh_counter[5] .power_up = "low";

cycloneive_lcell_comb \Add0~12 (
	.dataa(\refresh_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~5 (
	.dataa(\Add0~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~5_combout ),
	.cout());
defparam \refresh_counter~5 .lut_mask = 16'hAAFF;
defparam \refresh_counter~5 .sum_lutc_input = "datac";

dffeas \refresh_counter[6] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[6]~q ),
	.prn(vcc));
defparam \refresh_counter[6] .is_wysiwyg = "true";
defparam \refresh_counter[6] .power_up = "low";

cycloneive_lcell_comb \Add0~14 (
	.dataa(\refresh_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

dffeas \refresh_counter[7] (
	.clk(wire_pll7_clk_0),
	.d(\Add0~14_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[7]~q ),
	.prn(vcc));
defparam \refresh_counter[7] .is_wysiwyg = "true";
defparam \refresh_counter[7] .power_up = "low";

cycloneive_lcell_comb \Add0~16 (
	.dataa(\refresh_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'h5A5F;
defparam \Add0~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter[8]~13 (
	.dataa(\Add0~16_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\refresh_counter[8]~13_combout ),
	.cout());
defparam \refresh_counter[8]~13 .lut_mask = 16'h5555;
defparam \refresh_counter[8]~13 .sum_lutc_input = "datac";

dffeas \refresh_counter[8] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter[8]~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[8]~q ),
	.prn(vcc));
defparam \refresh_counter[8] .is_wysiwyg = "true";
defparam \refresh_counter[8] .power_up = "low";

cycloneive_lcell_comb \Add0~18 (
	.dataa(\refresh_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'h5AAF;
defparam \Add0~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~4 (
	.dataa(\Add0~18_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~4_combout ),
	.cout());
defparam \refresh_counter~4 .lut_mask = 16'hFF55;
defparam \refresh_counter~4 .sum_lutc_input = "datac";

dffeas \refresh_counter[9] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[9]~q ),
	.prn(vcc));
defparam \refresh_counter[9] .is_wysiwyg = "true";
defparam \refresh_counter[9] .power_up = "low";

cycloneive_lcell_comb \Add0~20 (
	.dataa(\refresh_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h5A5F;
defparam \Add0~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~1 (
	.dataa(\Add0~20_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~1_combout ),
	.cout());
defparam \refresh_counter~1 .lut_mask = 16'hFF55;
defparam \refresh_counter~1 .sum_lutc_input = "datac";

dffeas \refresh_counter[10] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[10]~q ),
	.prn(vcc));
defparam \refresh_counter[10] .is_wysiwyg = "true";
defparam \refresh_counter[10] .power_up = "low";

cycloneive_lcell_comb \Add0~22 (
	.dataa(\refresh_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~3 (
	.dataa(\Add0~22_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~3_combout ),
	.cout());
defparam \refresh_counter~3 .lut_mask = 16'hAAFF;
defparam \refresh_counter~3 .sum_lutc_input = "datac";

dffeas \refresh_counter[11] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[11]~q ),
	.prn(vcc));
defparam \refresh_counter[11] .is_wysiwyg = "true";
defparam \refresh_counter[11] .power_up = "low";

cycloneive_lcell_comb \Add0~24 (
	.dataa(\refresh_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'h5AAF;
defparam \Add0~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~2 (
	.dataa(\Add0~24_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~2_combout ),
	.cout());
defparam \refresh_counter~2 .lut_mask = 16'hAAFF;
defparam \refresh_counter~2 .sum_lutc_input = "datac";

dffeas \refresh_counter[12] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[12]~q ),
	.prn(vcc));
defparam \refresh_counter[12] .is_wysiwyg = "true";
defparam \refresh_counter[12] .power_up = "low";

cycloneive_lcell_comb \Add0~26 (
	.dataa(\refresh_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout());
defparam \Add0~26 .lut_mask = 16'h5A5A;
defparam \Add0~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \refresh_counter~0 (
	.dataa(\Add0~26_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~4_combout ),
	.cin(gnd),
	.combout(\refresh_counter~0_combout ),
	.cout());
defparam \refresh_counter~0 .lut_mask = 16'hFF55;
defparam \refresh_counter~0 .sum_lutc_input = "datac";

dffeas \refresh_counter[13] (
	.clk(wire_pll7_clk_0),
	.d(\refresh_counter~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_counter[13]~q ),
	.prn(vcc));
defparam \refresh_counter[13] .is_wysiwyg = "true";
defparam \refresh_counter[13] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\refresh_counter[13]~q ),
	.datab(\refresh_counter[10]~q ),
	.datac(\refresh_counter[12]~q ),
	.datad(\refresh_counter[11]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\refresh_counter[9]~q ),
	.datab(\refresh_counter[8]~q ),
	.datac(\refresh_counter[7]~q ),
	.datad(\refresh_counter[6]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\refresh_counter[4]~q ),
	.datab(\refresh_counter[5]~q ),
	.datac(\refresh_counter[3]~q ),
	.datad(\refresh_counter[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hBFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\refresh_counter[1]~q ),
	.datad(\refresh_counter[0]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h0FFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hFFFE;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_next.000~0 (
	.dataa(\i_next.000~q ),
	.datab(\i_state.000~q ),
	.datac(\i_state.101~q ),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\i_next.000~0_combout ),
	.cout());
defparam \i_next.000~0 .lut_mask = 16'hEFFF;
defparam \i_next.000~0 .sum_lutc_input = "datac";

dffeas \i_next.000 (
	.clk(wire_pll7_clk_0),
	.d(\i_next.000~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.000~q ),
	.prn(vcc));
defparam \i_next.000 .is_wysiwyg = "true";
defparam \i_next.000 .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\i_count[0]~0_combout ),
	.datab(\i_state.000~q ),
	.datac(\Equal0~4_combout ),
	.datad(\i_next.000~q ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFFFD;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \i_state.000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.000~q ),
	.prn(vcc));
defparam \i_state.000 .is_wysiwyg = "true";
defparam \i_state.000 .power_up = "low";

cycloneive_lcell_comb \Selector18~0 (
	.dataa(\i_next.111~q ),
	.datab(\i_state.101~q ),
	.datac(\i_state.011~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
defparam \Selector18~0 .lut_mask = 16'hFEFF;
defparam \Selector18~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hAAFF;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \i_state.001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.001~q ),
	.prn(vcc));
defparam \i_state.001 .is_wysiwyg = "true";
defparam \i_state.001 .power_up = "low";

cycloneive_lcell_comb \Selector16~0 (
	.dataa(\i_next.010~q ),
	.datab(\i_state.101~q ),
	.datac(\i_state.011~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
defparam \Selector16~0 .lut_mask = 16'hFEFF;
defparam \Selector16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(\i_state.010~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hAFFA;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas \i_refs[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(altera_reset_synchronizer_int_chain_out),
	.q(\i_refs[0]~q ),
	.prn(vcc));
defparam \i_refs[0] .is_wysiwyg = "true";
defparam \i_refs[0] .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\i_state.000~q ),
	.datab(\i_state.010~q ),
	.datac(\i_refs[1]~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEBBE;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \i_refs[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(altera_reset_synchronizer_int_chain_out),
	.q(\i_refs[1]~q ),
	.prn(vcc));
defparam \i_refs[1] .is_wysiwyg = "true";
defparam \i_refs[1] .power_up = "low";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\i_state.010~q ),
	.datab(\i_refs[2]~q ),
	.datac(\i_refs[1]~q ),
	.datad(\i_refs[0]~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEBBE;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(\Selector4~0_combout ),
	.datab(\i_state.000~q ),
	.datac(\i_refs[2]~q ),
	.datad(\i_state.010~q ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hFEFF;
defparam \Selector4~1 .sum_lutc_input = "datac";

dffeas \i_refs[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(altera_reset_synchronizer_int_chain_out),
	.q(\i_refs[2]~q ),
	.prn(vcc));
defparam \i_refs[2] .is_wysiwyg = "true";
defparam \i_refs[2] .power_up = "low";

cycloneive_lcell_comb \Selector18~1 (
	.dataa(\i_refs[0]~q ),
	.datab(gnd),
	.datac(\i_refs[2]~q ),
	.datad(\i_refs[1]~q ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
defparam \Selector18~1 .lut_mask = 16'hAFFF;
defparam \Selector18~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector16~1 (
	.dataa(\i_state.001~q ),
	.datab(\Selector16~0_combout ),
	.datac(\i_state.010~q ),
	.datad(\Selector18~1_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
defparam \Selector16~1 .lut_mask = 16'hFEFF;
defparam \Selector16~1 .sum_lutc_input = "datac";

dffeas \i_next.010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector16~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.010~q ),
	.prn(vcc));
defparam \i_next.010 .is_wysiwyg = "true";
defparam \i_next.010 .power_up = "low";

cycloneive_lcell_comb \i_count[0]~4 (
	.dataa(\i_state.010~q ),
	.datab(gnd),
	.datac(\i_state.011~q ),
	.datad(\i_count[0]~q ),
	.cin(gnd),
	.combout(\i_count[0]~4_combout ),
	.cout());
defparam \i_count[0]~4 .lut_mask = 16'hA0AF;
defparam \i_count[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_count[0]~1 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.101~q ),
	.cin(gnd),
	.combout(\i_count[0]~1_combout ),
	.cout());
defparam \i_count[0]~1 .lut_mask = 16'hAAFF;
defparam \i_count[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_count[0]~5 (
	.dataa(\i_count[0]~q ),
	.datab(\i_count[0]~4_combout ),
	.datac(\i_count[0]~1_combout ),
	.datad(\i_count[0]~0_combout ),
	.cin(gnd),
	.combout(\i_count[0]~5_combout ),
	.cout());
defparam \i_count[0]~5 .lut_mask = 16'hEFFE;
defparam \i_count[0]~5 .sum_lutc_input = "datac";

dffeas \i_count[0] (
	.clk(wire_pll7_clk_0),
	.d(\i_count[0]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[0]~q ),
	.prn(vcc));
defparam \i_count[0] .is_wysiwyg = "true";
defparam \i_count[0] .power_up = "low";

cycloneive_lcell_comb \i_count[1]~2 (
	.dataa(\i_count[1]~q ),
	.datab(\i_count[0]~q ),
	.datac(\i_state.010~q ),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\i_count[1]~2_combout ),
	.cout());
defparam \i_count[1]~2 .lut_mask = 16'hF9F6;
defparam \i_count[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_count[1]~3 (
	.dataa(\i_count[1]~q ),
	.datab(\i_count[1]~2_combout ),
	.datac(\i_count[0]~1_combout ),
	.datad(\i_count[0]~0_combout ),
	.cin(gnd),
	.combout(\i_count[1]~3_combout ),
	.cout());
defparam \i_count[1]~3 .lut_mask = 16'hEFFE;
defparam \i_count[1]~3 .sum_lutc_input = "datac";

dffeas \i_count[1] (
	.clk(wire_pll7_clk_0),
	.d(\i_count[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[1]~q ),
	.prn(vcc));
defparam \i_count[1] .is_wysiwyg = "true";
defparam \i_count[1] .power_up = "low";

cycloneive_lcell_comb \Selector13~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_count[1]~q ),
	.datac(\i_count[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hFEFE;
defparam \Selector13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector13~1 (
	.dataa(\i_state.111~q ),
	.datab(\i_count[2]~q ),
	.datac(\Selector13~0_combout ),
	.datad(\i_count[0]~1_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
defparam \Selector13~1 .lut_mask = 16'hFEFF;
defparam \Selector13~1 .sum_lutc_input = "datac";

dffeas \i_count[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector13~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_count[2]~q ),
	.prn(vcc));
defparam \i_count[2] .is_wysiwyg = "true";
defparam \i_count[2] .power_up = "low";

cycloneive_lcell_comb \Selector9~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_next.010~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hEFFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

dffeas \i_state.010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.010~q ),
	.prn(vcc));
defparam \i_state.010 .is_wysiwyg = "true";
defparam \i_state.010 .power_up = "low";

cycloneive_lcell_comb \Selector18~2 (
	.dataa(\Selector18~0_combout ),
	.datab(\i_state.010~q ),
	.datac(\Selector18~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
defparam \Selector18~2 .lut_mask = 16'hFEFE;
defparam \Selector18~2 .sum_lutc_input = "datac";

dffeas \i_next.111 (
	.clk(wire_pll7_clk_0),
	.d(\Selector18~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.111~q ),
	.prn(vcc));
defparam \i_next.111 .is_wysiwyg = "true";
defparam \i_next.111 .power_up = "low";

cycloneive_lcell_comb \Selector12~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_next.111~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'hEFFF;
defparam \Selector12~0 .sum_lutc_input = "datac";

dffeas \i_state.111 (
	.clk(wire_pll7_clk_0),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.111~q ),
	.prn(vcc));
defparam \i_state.111 .is_wysiwyg = "true";
defparam \i_state.111 .power_up = "low";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(\i_state.001~q ),
	.datab(\i_state.011~q ),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFFFE;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~1 (
	.dataa(\i_state.111~q ),
	.datab(\i_state.010~q ),
	.datac(\Selector10~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hFEFE;
defparam \Selector10~1 .sum_lutc_input = "datac";

dffeas \i_state.011 (
	.clk(wire_pll7_clk_0),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.011~q ),
	.prn(vcc));
defparam \i_state.011 .is_wysiwyg = "true";
defparam \i_state.011 .power_up = "low";

cycloneive_lcell_comb \i_count[0]~0 (
	.dataa(\i_state.011~q ),
	.datab(gnd),
	.datac(\i_count[2]~q ),
	.datad(\i_count[1]~q ),
	.cin(gnd),
	.combout(\i_count[0]~0_combout ),
	.cout());
defparam \i_count[0]~0 .lut_mask = 16'hAFFF;
defparam \i_count[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr6~0 (
	.dataa(\i_state.000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\i_state.011~q ),
	.cin(gnd),
	.combout(\WideOr6~0_combout ),
	.cout());
defparam \WideOr6~0 .lut_mask = 16'hAAFF;
defparam \WideOr6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector17~0 (
	.dataa(\i_state.111~q ),
	.datab(\i_next.101~q ),
	.datac(\i_state.101~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
defparam \Selector17~0 .lut_mask = 16'hFEFF;
defparam \Selector17~0 .sum_lutc_input = "datac";

dffeas \i_next.101 (
	.clk(wire_pll7_clk_0),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_next.101~q ),
	.prn(vcc));
defparam \i_next.101 .is_wysiwyg = "true";
defparam \i_next.101 .power_up = "low";

cycloneive_lcell_comb \i_state.101~0 (
	.dataa(\i_state.101~q ),
	.datab(\i_count[0]~0_combout ),
	.datac(\i_next.101~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\i_state.101~0_combout ),
	.cout());
defparam \i_state.101~0 .lut_mask = 16'hFEFE;
defparam \i_state.101~0 .sum_lutc_input = "datac";

dffeas \i_state.101 (
	.clk(wire_pll7_clk_0),
	.d(\i_state.101~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_state.101~q ),
	.prn(vcc));
defparam \i_state.101 .is_wysiwyg = "true";
defparam \i_state.101 .power_up = "low";

cycloneive_lcell_comb \init_done~0 (
	.dataa(\init_done~q ),
	.datab(\i_state.101~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\init_done~0_combout ),
	.cout());
defparam \init_done~0 .lut_mask = 16'hEEEE;
defparam \init_done~0 .sum_lutc_input = "datac";

dffeas init_done(
	.clk(wire_pll7_clk_0),
	.d(\init_done~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\init_done~q ),
	.prn(vcc));
defparam init_done.is_wysiwyg = "true";
defparam init_done.power_up = "low";

cycloneive_lcell_comb \Selector24~1 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\refresh_request~q ),
	.datad(\init_done~q ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
defparam \Selector24~1 .lut_mask = 16'h7FFF;
defparam \Selector24~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~0 (
	.dataa(\m_state.100000000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector32~0_combout ),
	.cout());
defparam \Selector32~0 .lut_mask = 16'hAAFF;
defparam \Selector32~0 .sum_lutc_input = "datac";

dffeas active_rnw(
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_rnw~q ),
	.prn(vcc));
defparam active_rnw.is_wysiwyg = "true";
defparam active_rnw.power_up = "low";

cycloneive_lcell_comb \Selector25~5 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(gnd),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
defparam \Selector25~5 .lut_mask = 16'hEEFF;
defparam \Selector25~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector25~6 (
	.dataa(\init_done~q ),
	.datab(\m_state.000000001~q ),
	.datac(\Selector25~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector25~6_combout ),
	.cout());
defparam \Selector25~6 .lut_mask = 16'hFBFB;
defparam \Selector25~6 .sum_lutc_input = "datac";

dffeas \m_state.000000010 (
	.clk(wire_pll7_clk_0),
	.d(\Selector25~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000010~q ),
	.prn(vcc));
defparam \m_state.000000010 .is_wysiwyg = "true";
defparam \m_state.000000010 .power_up = "low";

dffeas \active_addr[10] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[10]~q ),
	.prn(vcc));
defparam \active_addr[10] .is_wysiwyg = "true";
defparam \active_addr[10] .power_up = "low";

cycloneive_lcell_comb \pending~0 (
	.dataa(\active_rnw~q ),
	.datab(\active_addr[10]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.cin(gnd),
	.combout(\pending~0_combout ),
	.cout());
defparam \pending~0 .lut_mask = 16'h6996;
defparam \pending~0 .sum_lutc_input = "datac";

dffeas \active_addr[24] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[24]~q ),
	.prn(vcc));
defparam \active_addr[24] .is_wysiwyg = "true";
defparam \active_addr[24] .power_up = "low";

cycloneive_lcell_comb \pending~1 (
	.dataa(\active_addr[11]~q ),
	.datab(\active_addr[24]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[47]~3_combout ),
	.cin(gnd),
	.combout(\pending~1_combout ),
	.cout());
defparam \pending~1 .lut_mask = 16'h6996;
defparam \pending~1 .sum_lutc_input = "datac";

dffeas \active_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[48]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[12]~q ),
	.prn(vcc));
defparam \active_addr[12] .is_wysiwyg = "true";
defparam \active_addr[12] .power_up = "low";

dffeas \active_addr[13] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[49]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[13]~q ),
	.prn(vcc));
defparam \active_addr[13] .is_wysiwyg = "true";
defparam \active_addr[13] .power_up = "low";

cycloneive_lcell_comb \pending~2 (
	.dataa(\active_addr[12]~q ),
	.datab(\active_addr[13]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[49]~4_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[48]~5_combout ),
	.cin(gnd),
	.combout(\pending~2_combout ),
	.cout());
defparam \pending~2 .lut_mask = 16'h6996;
defparam \pending~2 .sum_lutc_input = "datac";

dffeas \active_addr[14] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[50]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[14]~q ),
	.prn(vcc));
defparam \active_addr[14] .is_wysiwyg = "true";
defparam \active_addr[14] .power_up = "low";

dffeas \active_addr[15] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[51]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[15]~q ),
	.prn(vcc));
defparam \active_addr[15] .is_wysiwyg = "true";
defparam \active_addr[15] .power_up = "low";

cycloneive_lcell_comb \pending~3 (
	.dataa(\active_addr[14]~q ),
	.datab(\active_addr[15]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[51]~6_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[50]~7_combout ),
	.cin(gnd),
	.combout(\pending~3_combout ),
	.cout());
defparam \pending~3 .lut_mask = 16'h6996;
defparam \pending~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~4 (
	.dataa(\pending~0_combout ),
	.datab(\pending~1_combout ),
	.datac(\pending~2_combout ),
	.datad(\pending~3_combout ),
	.cin(gnd),
	.combout(\pending~4_combout ),
	.cout());
defparam \pending~4 .lut_mask = 16'hFFFE;
defparam \pending~4 .sum_lutc_input = "datac";

dffeas \active_addr[16] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[52]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[16]~q ),
	.prn(vcc));
defparam \active_addr[16] .is_wysiwyg = "true";
defparam \active_addr[16] .power_up = "low";

dffeas \active_addr[17] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[53]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[17]~q ),
	.prn(vcc));
defparam \active_addr[17] .is_wysiwyg = "true";
defparam \active_addr[17] .power_up = "low";

cycloneive_lcell_comb \pending~5 (
	.dataa(\active_addr[16]~q ),
	.datab(\active_addr[17]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[53]~8_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[52]~9_combout ),
	.cin(gnd),
	.combout(\pending~5_combout ),
	.cout());
defparam \pending~5 .lut_mask = 16'h6996;
defparam \pending~5 .sum_lutc_input = "datac";

dffeas \active_addr[18] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[54]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[18]~q ),
	.prn(vcc));
defparam \active_addr[18] .is_wysiwyg = "true";
defparam \active_addr[18] .power_up = "low";

dffeas \active_addr[19] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[55]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[19]~q ),
	.prn(vcc));
defparam \active_addr[19] .is_wysiwyg = "true";
defparam \active_addr[19] .power_up = "low";

cycloneive_lcell_comb \pending~6 (
	.dataa(\active_addr[18]~q ),
	.datab(\active_addr[19]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[55]~10_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[54]~11_combout ),
	.cin(gnd),
	.combout(\pending~6_combout ),
	.cout());
defparam \pending~6 .lut_mask = 16'h6996;
defparam \pending~6 .sum_lutc_input = "datac";

dffeas \active_addr[20] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[56]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[20]~q ),
	.prn(vcc));
defparam \active_addr[20] .is_wysiwyg = "true";
defparam \active_addr[20] .power_up = "low";

dffeas \active_addr[21] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[57]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[21]~q ),
	.prn(vcc));
defparam \active_addr[21] .is_wysiwyg = "true";
defparam \active_addr[21] .power_up = "low";

cycloneive_lcell_comb \pending~7 (
	.dataa(\active_addr[20]~q ),
	.datab(\active_addr[21]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[57]~12_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[56]~13_combout ),
	.cin(gnd),
	.combout(\pending~7_combout ),
	.cout());
defparam \pending~7 .lut_mask = 16'h6996;
defparam \pending~7 .sum_lutc_input = "datac";

dffeas \active_addr[22] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[58]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[22]~q ),
	.prn(vcc));
defparam \active_addr[22] .is_wysiwyg = "true";
defparam \active_addr[22] .power_up = "low";

dffeas \active_addr[23] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[59]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[23]~q ),
	.prn(vcc));
defparam \active_addr[23] .is_wysiwyg = "true";
defparam \active_addr[23] .power_up = "low";

cycloneive_lcell_comb \pending~8 (
	.dataa(\active_addr[22]~q ),
	.datab(\active_addr[23]~q ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|rd_data[59]~14_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[58]~15_combout ),
	.cin(gnd),
	.combout(\pending~8_combout ),
	.cout());
defparam \pending~8 .lut_mask = 16'h6996;
defparam \pending~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~9 (
	.dataa(\pending~5_combout ),
	.datab(\pending~6_combout ),
	.datac(\pending~7_combout ),
	.datad(\pending~8_combout ),
	.cin(gnd),
	.combout(\pending~9_combout ),
	.cout());
defparam \pending~9 .lut_mask = 16'hFFFE;
defparam \pending~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_next~19 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\active_cs_n~q ),
	.datac(\pending~4_combout ),
	.datad(\pending~9_combout ),
	.cin(gnd),
	.combout(\m_next~19_combout ),
	.cout());
defparam \m_next~19 .lut_mask = 16'hEFFF;
defparam \m_next~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector25~4 (
	.dataa(\init_done~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
defparam \Selector25~4 .lut_mask = 16'hAAFF;
defparam \Selector25~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \pending~10 (
	.dataa(\pending~4_combout ),
	.datab(\pending~9_combout ),
	.datac(gnd),
	.datad(\active_cs_n~q ),
	.cin(gnd),
	.combout(\pending~10_combout ),
	.cout());
defparam \pending~10 .lut_mask = 16'hEEFF;
defparam \pending~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~0 (
	.dataa(\m_state.100000000~q ),
	.datab(\pending~10_combout ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hEFFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_next~20 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(\pending~10_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\m_next~20_combout ),
	.cout());
defparam \m_next~20 .lut_mask = 16'hFFFE;
defparam \m_next~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector29~0 (
	.dataa(\m_state.100000000~q ),
	.datab(\active_cs_n~q ),
	.datac(\pending~4_combout ),
	.datad(\pending~9_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
defparam \Selector29~0 .lut_mask = 16'hEFFF;
defparam \Selector29~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~0 (
	.dataa(\Selector24~0_combout ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\refresh_request~q ),
	.datad(\m_state.100000000~q ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
defparam \Selector27~0 .lut_mask = 16'hBFFF;
defparam \Selector27~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~0 (
	.dataa(\m_state.000000010~q ),
	.datab(\Selector34~0_combout ),
	.datac(gnd),
	.datad(\active_rnw~q ),
	.cin(gnd),
	.combout(\Selector35~0_combout ),
	.cout());
defparam \Selector35~0 .lut_mask = 16'hEEFF;
defparam \Selector35~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~2 (
	.dataa(\m_state.000000010~q ),
	.datab(\refresh_request~q ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector34~2_combout ),
	.cout());
defparam \Selector34~2 .lut_mask = 16'hEFFF;
defparam \Selector34~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~3 (
	.dataa(\Selector34~2_combout ),
	.datab(\m_next~20_combout ),
	.datac(\WideOr9~0_combout ),
	.datad(\Selector34~0_combout ),
	.cin(gnd),
	.combout(\Selector34~3_combout ),
	.cout());
defparam \Selector34~3 .lut_mask = 16'hEFFF;
defparam \Selector34~3 .sum_lutc_input = "datac";

dffeas \m_next.000010000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector35~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector34~3_combout ),
	.q(\m_next.000010000~q ),
	.prn(vcc));
defparam \m_next.000010000 .is_wysiwyg = "true";
defparam \m_next.000010000 .power_up = "low";

cycloneive_lcell_comb \Selector27~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\pending~10_combout ),
	.datac(\m_state.100000000~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
defparam \Selector27~1 .lut_mask = 16'hFEFF;
defparam \Selector27~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector28~0 (
	.dataa(\Selector27~0_combout ),
	.datab(\m_next.000010000~q ),
	.datac(\Selector27~1_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
defparam \Selector28~0 .lut_mask = 16'hFEFF;
defparam \Selector28~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~3 (
	.dataa(\refresh_request~q ),
	.datab(\pending~combout ),
	.datac(\m_state.000000001~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
defparam \Selector27~3 .lut_mask = 16'hFEFF;
defparam \Selector27~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~4 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datab(\refresh_request~q ),
	.datac(\init_done~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
defparam \Selector27~4 .lut_mask = 16'hEFFF;
defparam \Selector27~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr8~0 (
	.dataa(gnd),
	.datab(\m_state.000000010~q ),
	.datac(\m_state.001000000~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\WideOr8~0_combout ),
	.cout());
defparam \WideOr8~0 .lut_mask = 16'h3FFF;
defparam \WideOr8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~5 (
	.dataa(\m_state.100000000~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\refresh_request~q ),
	.datad(\WideOr8~0_combout ),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
defparam \Selector27~5 .lut_mask = 16'hFEFF;
defparam \Selector27~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~6 (
	.dataa(\Selector24~0_combout ),
	.datab(\Selector27~3_combout ),
	.datac(\Selector27~4_combout ),
	.datad(\Selector27~5_combout ),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
defparam \Selector27~6 .lut_mask = 16'hFFFE;
defparam \Selector27~6 .sum_lutc_input = "datac";

dffeas \m_state.000010000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector27~6_combout ),
	.q(\m_state.000010000~q ),
	.prn(vcc));
defparam \m_state.000010000 .is_wysiwyg = "true";
defparam \m_state.000010000 .power_up = "low";

cycloneive_lcell_comb \Selector39~0 (
	.dataa(\m_next~20_combout ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000001000~q ),
	.datad(\Selector38~0_combout ),
	.cin(gnd),
	.combout(\Selector39~0_combout ),
	.cout());
defparam \Selector39~0 .lut_mask = 16'hBFFF;
defparam \Selector39~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~1 (
	.dataa(\m_count[1]~q ),
	.datab(\m_state.000000100~q ),
	.datac(\m_state.000100000~q ),
	.datad(\m_count[0]~q ),
	.cin(gnd),
	.combout(\Selector39~1_combout ),
	.cout());
defparam \Selector39~1 .lut_mask = 16'hBFFF;
defparam \Selector39~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~2 (
	.dataa(\m_state.000000001~q ),
	.datab(\Selector39~0_combout ),
	.datac(\Selector39~1_combout ),
	.datad(\m_state.001000000~q ),
	.cin(gnd),
	.combout(\Selector39~2_combout ),
	.cout());
defparam \Selector39~2 .lut_mask = 16'hFEFF;
defparam \Selector39~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~3 (
	.dataa(\m_count[0]~q ),
	.datab(\m_state.000000001~q ),
	.datac(\init_done~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector39~3_combout ),
	.cout());
defparam \Selector39~3 .lut_mask = 16'hEFFF;
defparam \Selector39~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~4 (
	.dataa(\Selector39~3_combout ),
	.datab(\m_state.000000100~q ),
	.datac(\m_count[1]~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector39~4_combout ),
	.cout());
defparam \Selector39~4 .lut_mask = 16'hBFFF;
defparam \Selector39~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector39~5 (
	.dataa(\Selector39~2_combout ),
	.datab(\Selector39~4_combout ),
	.datac(\m_state.000001000~q ),
	.datad(\m_next~20_combout ),
	.cin(gnd),
	.combout(\Selector39~5_combout ),
	.cout());
defparam \Selector39~5 .lut_mask = 16'hEFFF;
defparam \Selector39~5 .sum_lutc_input = "datac";

dffeas \m_count[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector39~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[0]~q ),
	.prn(vcc));
defparam \m_count[0] .is_wysiwyg = "true";
defparam \m_count[0] .power_up = "low";

cycloneive_lcell_comb \Selector38~1 (
	.dataa(\m_count[1]~q ),
	.datab(\m_count[0]~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector38~1_combout ),
	.cout());
defparam \Selector38~1 .lut_mask = 16'hFFFE;
defparam \Selector38~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~2 (
	.dataa(\m_state.010000000~q ),
	.datab(\Selector38~1_combout ),
	.datac(\m_state.000001000~q ),
	.datad(\m_next~20_combout ),
	.cin(gnd),
	.combout(\Selector38~2_combout ),
	.cout());
defparam \Selector38~2 .lut_mask = 16'hFFFE;
defparam \Selector38~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~3 (
	.dataa(\m_state.001000000~q ),
	.datab(\init_done~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector38~3_combout ),
	.cout());
defparam \Selector38~3 .lut_mask = 16'hBFFF;
defparam \Selector38~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector38~4 (
	.dataa(\Selector38~2_combout ),
	.datab(\m_count[1]~q ),
	.datac(\Selector38~3_combout ),
	.datad(\Selector39~0_combout ),
	.cin(gnd),
	.combout(\Selector38~4_combout ),
	.cout());
defparam \Selector38~4 .lut_mask = 16'hFEFF;
defparam \Selector38~4 .sum_lutc_input = "datac";

dffeas \m_count[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector38~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_count[1]~q ),
	.prn(vcc));
defparam \m_count[1] .is_wysiwyg = "true";
defparam \m_count[1] .power_up = "low";

cycloneive_lcell_comb \Selector29~1 (
	.dataa(\m_state.000100000~q ),
	.datab(\Selector29~0_combout ),
	.datac(\Selector25~5_combout ),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
defparam \Selector29~1 .lut_mask = 16'hFFFE;
defparam \Selector29~1 .sum_lutc_input = "datac";

dffeas \m_state.000100000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector29~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000100000~q ),
	.prn(vcc));
defparam \m_state.000100000 .is_wysiwyg = "true";
defparam \m_state.000100000 .power_up = "low";

cycloneive_lcell_comb \Selector30~0 (
	.dataa(\m_state.000100000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
defparam \Selector30~0 .lut_mask = 16'hAAFF;
defparam \Selector30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector30~1 (
	.dataa(\Selector30~0_combout ),
	.datab(\init_done~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector30~1_combout ),
	.cout());
defparam \Selector30~1 .lut_mask = 16'hFEFF;
defparam \Selector30~1 .sum_lutc_input = "datac";

dffeas \m_state.001000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector30~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.001000000~q ),
	.prn(vcc));
defparam \m_state.001000000 .is_wysiwyg = "true";
defparam \m_state.001000000 .power_up = "low";

cycloneive_lcell_comb \Selector33~0 (
	.dataa(gnd),
	.datab(\m_state.001000000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\Selector33~0_combout ),
	.cout());
defparam \Selector33~0 .lut_mask = 16'h3FFF;
defparam \Selector33~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~0 (
	.dataa(\Selector38~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\m_next~20_combout ),
	.datad(\Selector33~0_combout ),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
defparam \Selector36~0 .lut_mask = 16'hBFFF;
defparam \Selector36~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~1 (
	.dataa(\Selector25~4_combout ),
	.datab(\m_next.010000000~q ),
	.datac(\Selector36~0_combout ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector36~1_combout ),
	.cout());
defparam \Selector36~1 .lut_mask = 16'hFFFE;
defparam \Selector36~1 .sum_lutc_input = "datac";

dffeas \m_next.010000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector36~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.010000000~q ),
	.prn(vcc));
defparam \m_next.010000000 .is_wysiwyg = "true";
defparam \m_next.010000000 .power_up = "low";

cycloneive_lcell_comb \Selector31~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_next.010000000~q ),
	.datac(gnd),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
defparam \Selector31~0 .lut_mask = 16'hEEFF;
defparam \Selector31~0 .sum_lutc_input = "datac";

dffeas \m_state.010000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.010000000~q ),
	.prn(vcc));
defparam \m_state.010000000 .is_wysiwyg = "true";
defparam \m_state.010000000 .power_up = "low";

cycloneive_lcell_comb \Selector34~0 (
	.dataa(\refresh_request~q ),
	.datab(\m_next~19_combout ),
	.datac(\m_state.100000000~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector34~0_combout ),
	.cout());
defparam \Selector34~0 .lut_mask = 16'h7FFF;
defparam \Selector34~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector34~1 (
	.dataa(\active_rnw~q ),
	.datab(\m_state.000000010~q ),
	.datac(\Selector34~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector34~1_combout ),
	.cout());
defparam \Selector34~1 .lut_mask = 16'hFEFE;
defparam \Selector34~1 .sum_lutc_input = "datac";

dffeas \m_next.000001000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector34~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector34~3_combout ),
	.q(\m_next.000001000~q ),
	.prn(vcc));
defparam \m_next.000001000 .is_wysiwyg = "true";
defparam \m_next.000001000 .power_up = "low";

cycloneive_lcell_comb \Selector27~2 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[61]~1_combout ),
	.datab(\m_next.000001000~q ),
	.datac(\Selector27~0_combout ),
	.datad(\Selector27~1_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
defparam \Selector27~2 .lut_mask = 16'hFFFE;
defparam \Selector27~2 .sum_lutc_input = "datac";

dffeas \m_state.000001000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector27~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector27~6_combout ),
	.q(\m_state.000001000~q ),
	.prn(vcc));
defparam \m_state.000001000 .is_wysiwyg = "true";
defparam \m_state.000001000 .power_up = "low";

cycloneive_lcell_comb \WideOr9~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\m_state.000001000~q ),
	.datad(\m_state.000010000~q ),
	.cin(gnd),
	.combout(\WideOr9~0_combout ),
	.cout());
defparam \WideOr9~0 .lut_mask = 16'h0FFF;
defparam \WideOr9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~1 (
	.dataa(\Selector32~0_combout ),
	.datab(\pending~combout ),
	.datac(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector32~1_combout ),
	.cout());
defparam \Selector32~1 .lut_mask = 16'hEFFF;
defparam \Selector32~1 .sum_lutc_input = "datac";

dffeas \m_state.100000000 (
	.clk(wire_pll7_clk_0),
	.d(\Selector32~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.100000000~q ),
	.prn(vcc));
defparam \m_state.100000000 .is_wysiwyg = "true";
defparam \m_state.100000000 .power_up = "low";

cycloneive_lcell_comb \Selector26~0 (
	.dataa(\m_state.000000100~q ),
	.datab(\m_state.100000000~q ),
	.datac(\refresh_request~q ),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
defparam \Selector26~0 .lut_mask = 16'hFFFE;
defparam \Selector26~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~1 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
defparam \Selector26~1 .lut_mask = 16'hFFFE;
defparam \Selector26~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector26~2 (
	.dataa(\Selector26~0_combout ),
	.datab(\Selector26~1_combout ),
	.datac(\pending~combout ),
	.datad(\WideOr8~0_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
defparam \Selector26~2 .lut_mask = 16'hEFFF;
defparam \Selector26~2 .sum_lutc_input = "datac";

dffeas \m_state.000000100 (
	.clk(wire_pll7_clk_0),
	.d(\Selector26~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000100~q ),
	.prn(vcc));
defparam \m_state.000000100 .is_wysiwyg = "true";
defparam \m_state.000000100 .power_up = "low";

cycloneive_lcell_comb \Selector24~0 (
	.dataa(\m_state.000000100~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\m_count[1]~q ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
defparam \Selector24~0 .lut_mask = 16'hAAFF;
defparam \Selector24~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~1 (
	.dataa(\m_state.001000000~q ),
	.datab(\m_state.000000100~q ),
	.datac(\m_state.000100000~q ),
	.datad(\m_state.100000000~q ),
	.cin(gnd),
	.combout(\Selector33~1_combout ),
	.cout());
defparam \Selector33~1 .lut_mask = 16'hFFFE;
defparam \Selector33~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~2 (
	.dataa(\Selector33~1_combout ),
	.datab(\m_state.000000001~q ),
	.datac(\refresh_request~q ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector33~2_combout ),
	.cout());
defparam \Selector33~2 .lut_mask = 16'hBFFF;
defparam \Selector33~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~3 (
	.dataa(\Selector33~2_combout ),
	.datab(\init_done~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_next.000000001~q ),
	.cin(gnd),
	.combout(\Selector33~3_combout ),
	.cout());
defparam \Selector33~3 .lut_mask = 16'hBFFF;
defparam \Selector33~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~4 (
	.dataa(\Selector33~3_combout ),
	.datab(\m_next~20_combout ),
	.datac(\WideOr9~0_combout ),
	.datad(\Selector34~0_combout ),
	.cin(gnd),
	.combout(\Selector33~4_combout ),
	.cout());
defparam \Selector33~4 .lut_mask = 16'hFFF7;
defparam \Selector33~4 .sum_lutc_input = "datac";

dffeas \m_next.000000001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector33~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_next.000000001~q ),
	.prn(vcc));
defparam \m_next.000000001 .is_wysiwyg = "true";
defparam \m_next.000000001 .power_up = "low";

cycloneive_lcell_comb \Selector24~2 (
	.dataa(\Selector24~1_combout ),
	.datab(\Selector24~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\m_next.000000001~q ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
defparam \Selector24~2 .lut_mask = 16'hFFF7;
defparam \Selector24~2 .sum_lutc_input = "datac";

dffeas \m_state.000000001 (
	.clk(wire_pll7_clk_0),
	.d(\Selector24~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_state.000000001~q ),
	.prn(vcc));
defparam \m_state.000000001 .is_wysiwyg = "true";
defparam \m_state.000000001 .power_up = "low";

cycloneive_lcell_comb \Selector23~0 (
	.dataa(\m_state.000000001~q ),
	.datab(\ack_refresh_request~q ),
	.datac(\m_state.010000000~q ),
	.datad(\init_done~q ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
defparam \Selector23~0 .lut_mask = 16'hFEFF;
defparam \Selector23~0 .sum_lutc_input = "datac";

dffeas ack_refresh_request(
	.clk(wire_pll7_clk_0),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ack_refresh_request~q ),
	.prn(vcc));
defparam ack_refresh_request.is_wysiwyg = "true";
defparam ack_refresh_request.power_up = "low";

cycloneive_lcell_comb \refresh_request~0 (
	.dataa(\init_done~q ),
	.datab(\refresh_request~q ),
	.datac(\Equal0~4_combout ),
	.datad(\ack_refresh_request~q ),
	.cin(gnd),
	.combout(\refresh_request~0_combout ),
	.cout());
defparam \refresh_request~0 .lut_mask = 16'hFEFF;
defparam \refresh_request~0 .sum_lutc_input = "datac";

dffeas refresh_request(
	.clk(wire_pll7_clk_0),
	.d(\refresh_request~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_request~q ),
	.prn(vcc));
defparam refresh_request.is_wysiwyg = "true";
defparam refresh_request.power_up = "low";

cycloneive_lcell_comb \active_cs_n~0 (
	.dataa(altera_reset_synchronizer_int_chain_out),
	.datab(\init_done~q ),
	.datac(gnd),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\active_cs_n~0_combout ),
	.cout());
defparam \active_cs_n~0 .lut_mask = 16'hEEFF;
defparam \active_cs_n~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_cs_n~1 (
	.dataa(\refresh_request~q ),
	.datab(\active_cs_n~q ),
	.datac(\active_cs_n~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.cin(gnd),
	.combout(\active_cs_n~1_combout ),
	.cout());
defparam \active_cs_n~1 .lut_mask = 16'hACFF;
defparam \active_cs_n~1 .sum_lutc_input = "datac";

dffeas active_cs_n(
	.clk(wire_pll7_clk_0),
	.d(\active_cs_n~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\active_cs_n~q ),
	.prn(vcc));
defparam active_cs_n.is_wysiwyg = "true";
defparam active_cs_n.power_up = "low";

cycloneive_lcell_comb pending(
	.dataa(\active_cs_n~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|Equal1~0_combout ),
	.datac(\pending~4_combout ),
	.datad(\pending~9_combout ),
	.cin(gnd),
	.combout(\pending~combout ),
	.cout());
defparam pending.lut_mask = 16'hBFFF;
defparam pending.sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~2 (
	.dataa(\pending~combout ),
	.datab(\refresh_request~q ),
	.datac(\m_state.000001000~q ),
	.datad(\m_state.000010000~q ),
	.cin(gnd),
	.combout(\active_rnw~2_combout ),
	.cout());
defparam \active_rnw~2 .lut_mask = 16'hEFFF;
defparam \active_rnw~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~4 (
	.dataa(\init_done~q ),
	.datab(\m_state.000000001~q ),
	.datac(\m_state.100000000~q ),
	.datad(\Selector25~5_combout ),
	.cin(gnd),
	.combout(\active_rnw~4_combout ),
	.cout());
defparam \active_rnw~4 .lut_mask = 16'hDFFF;
defparam \active_rnw~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \active_rnw~3 (
	.dataa(\active_rnw~2_combout ),
	.datab(\Selector29~0_combout ),
	.datac(\active_rnw~4_combout ),
	.datad(altera_reset_synchronizer_int_chain_out),
	.cin(gnd),
	.combout(\active_rnw~3_combout ),
	.cout());
defparam \active_rnw~3 .lut_mask = 16'hFF7F;
defparam \active_rnw~3 .sum_lutc_input = "datac";

dffeas \active_addr[11] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[47]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[11]~q ),
	.prn(vcc));
defparam \active_addr[11] .is_wysiwyg = "true";
defparam \active_addr[11] .power_up = "low";

cycloneive_lcell_comb \Selector41~0 (
	.dataa(\m_state.100000000~q ),
	.datab(entries_1),
	.datac(entries_0),
	.datad(\refresh_request~q ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
defparam \Selector41~0 .lut_mask = 16'hFEFF;
defparam \Selector41~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector41~1 (
	.dataa(\Selector25~6_combout ),
	.datab(\pending~10_combout ),
	.datac(\Selector41~0_combout ),
	.datad(\active_rnw~2_combout ),
	.cin(gnd),
	.combout(\Selector41~1_combout ),
	.cout());
defparam \Selector41~1 .lut_mask = 16'hFEFF;
defparam \Selector41~1 .sum_lutc_input = "datac";

dffeas f_pop(
	.clk(wire_pll7_clk_0),
	.d(\Selector41~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\f_pop~q ),
	.prn(vcc));
defparam f_pop.is_wysiwyg = "true";
defparam f_pop.power_up = "low";

cycloneive_lcell_comb \m_addr[3]~0 (
	.dataa(\m_state.000000010~q ),
	.datab(\WideOr9~0_combout ),
	.datac(\f_pop~q ),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\m_addr[3]~0_combout ),
	.cout());
defparam \m_addr[3]~0 .lut_mask = 16'hB8FF;
defparam \m_addr[3]~0 .sum_lutc_input = "datac";

dffeas \active_addr[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[36]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[0]~q ),
	.prn(vcc));
defparam \active_addr[0] .is_wysiwyg = "true";
defparam \active_addr[0] .power_up = "low";

dffeas \i_addr[12] (
	.clk(wire_pll7_clk_0),
	.d(\i_state.111~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_addr[12]~q ),
	.prn(vcc));
defparam \i_addr[12] .is_wysiwyg = "true";
defparam \i_addr[12] .power_up = "low";

cycloneive_lcell_comb \Selector116~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[0]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector116~0_combout ),
	.cout());
defparam \Selector116~0 .lut_mask = 16'hDEFF;
defparam \Selector116~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector116~1 (
	.dataa(\active_addr[11]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector116~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[36]~16_combout ),
	.cin(gnd),
	.combout(\Selector116~1_combout ),
	.cout());
defparam \Selector116~1 .lut_mask = 16'hFFBE;
defparam \Selector116~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_addr[3]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.000100000~q ),
	.cin(gnd),
	.combout(\m_addr[3]~1_combout ),
	.cout());
defparam \m_addr[3]~1 .lut_mask = 16'h0FFF;
defparam \m_addr[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_addr[3]~2 (
	.dataa(\m_state.010000000~q ),
	.datab(\m_state.100000000~q ),
	.datac(\Selector25~4_combout ),
	.datad(\m_addr[3]~1_combout ),
	.cin(gnd),
	.combout(\m_addr[3]~2_combout ),
	.cout());
defparam \m_addr[3]~2 .lut_mask = 16'hFF7F;
defparam \m_addr[3]~2 .sum_lutc_input = "datac";

dffeas \active_addr[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[37]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[1]~q ),
	.prn(vcc));
defparam \active_addr[1] .is_wysiwyg = "true";
defparam \active_addr[1] .power_up = "low";

cycloneive_lcell_comb \Selector115~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[1]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector115~0_combout ),
	.cout());
defparam \Selector115~0 .lut_mask = 16'hDEFF;
defparam \Selector115~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector115~1 (
	.dataa(\active_addr[12]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector115~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[37]~17_combout ),
	.cin(gnd),
	.combout(\Selector115~1_combout ),
	.cout());
defparam \Selector115~1 .lut_mask = 16'hFFBE;
defparam \Selector115~1 .sum_lutc_input = "datac";

dffeas \active_addr[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[38]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[2]~q ),
	.prn(vcc));
defparam \active_addr[2] .is_wysiwyg = "true";
defparam \active_addr[2] .power_up = "low";

cycloneive_lcell_comb \Selector114~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[2]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector114~0_combout ),
	.cout());
defparam \Selector114~0 .lut_mask = 16'hDEFF;
defparam \Selector114~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector114~1 (
	.dataa(\active_addr[13]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector114~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[38]~18_combout ),
	.cin(gnd),
	.combout(\Selector114~1_combout ),
	.cout());
defparam \Selector114~1 .lut_mask = 16'hFFBE;
defparam \Selector114~1 .sum_lutc_input = "datac";

dffeas \active_addr[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[39]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[3]~q ),
	.prn(vcc));
defparam \active_addr[3] .is_wysiwyg = "true";
defparam \active_addr[3] .power_up = "low";

cycloneive_lcell_comb \Selector113~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[3]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector113~0_combout ),
	.cout());
defparam \Selector113~0 .lut_mask = 16'hDEFF;
defparam \Selector113~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector113~1 (
	.dataa(\active_addr[14]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector113~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[39]~19_combout ),
	.cin(gnd),
	.combout(\Selector113~1_combout ),
	.cout());
defparam \Selector113~1 .lut_mask = 16'hFFBE;
defparam \Selector113~1 .sum_lutc_input = "datac";

dffeas \active_addr[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[40]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[4]~q ),
	.prn(vcc));
defparam \active_addr[4] .is_wysiwyg = "true";
defparam \active_addr[4] .power_up = "low";

cycloneive_lcell_comb \Selector112~0 (
	.dataa(\active_addr[4]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[40]~20_combout ),
	.datac(\f_pop~q ),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\Selector112~0_combout ),
	.cout());
defparam \Selector112~0 .lut_mask = 16'hEFFE;
defparam \Selector112~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector112~1 (
	.dataa(\active_addr[15]~q ),
	.datab(\Selector112~0_combout ),
	.datac(\WideOr9~0_combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector112~1_combout ),
	.cout());
defparam \Selector112~1 .lut_mask = 16'hACFF;
defparam \Selector112~1 .sum_lutc_input = "datac";

dffeas \active_addr[5] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[41]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[5]~q ),
	.prn(vcc));
defparam \active_addr[5] .is_wysiwyg = "true";
defparam \active_addr[5] .power_up = "low";

cycloneive_lcell_comb f_select(
	.dataa(\f_pop~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\f_select~combout ),
	.cout());
defparam f_select.lut_mask = 16'hAAFF;
defparam f_select.sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector111~0 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[41]~21_combout ),
	.datab(\active_addr[5]~q ),
	.datac(\f_select~combout ),
	.datad(\WideOr9~0_combout ),
	.cin(gnd),
	.combout(\Selector111~0_combout ),
	.cout());
defparam \Selector111~0 .lut_mask = 16'hACFF;
defparam \Selector111~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector111~1 (
	.dataa(\Selector111~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\active_addr[16]~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector111~1_combout ),
	.cout());
defparam \Selector111~1 .lut_mask = 16'hFEFF;
defparam \Selector111~1 .sum_lutc_input = "datac";

dffeas \active_addr[6] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[42]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[6]~q ),
	.prn(vcc));
defparam \active_addr[6] .is_wysiwyg = "true";
defparam \active_addr[6] .power_up = "low";

cycloneive_lcell_comb \Selector110~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[6]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector110~0_combout ),
	.cout());
defparam \Selector110~0 .lut_mask = 16'hDEFF;
defparam \Selector110~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector110~1 (
	.dataa(\active_addr[17]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector110~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[42]~22_combout ),
	.cin(gnd),
	.combout(\Selector110~1_combout ),
	.cout());
defparam \Selector110~1 .lut_mask = 16'hFFBE;
defparam \Selector110~1 .sum_lutc_input = "datac";

dffeas \active_addr[7] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[43]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[7]~q ),
	.prn(vcc));
defparam \active_addr[7] .is_wysiwyg = "true";
defparam \active_addr[7] .power_up = "low";

cycloneive_lcell_comb \Selector109~0 (
	.dataa(\WideOr9~0_combout ),
	.datab(\active_addr[18]~q ),
	.datac(\m_addr[3]~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector109~0_combout ),
	.cout());
defparam \Selector109~0 .lut_mask = 16'hDEFF;
defparam \Selector109~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector109~1 (
	.dataa(\active_addr[7]~q ),
	.datab(\WideOr9~0_combout ),
	.datac(\Selector109~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[43]~23_combout ),
	.cin(gnd),
	.combout(\Selector109~1_combout ),
	.cout());
defparam \Selector109~1 .lut_mask = 16'hFFBE;
defparam \Selector109~1 .sum_lutc_input = "datac";

dffeas \active_addr[8] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[44]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[8]~q ),
	.prn(vcc));
defparam \active_addr[8] .is_wysiwyg = "true";
defparam \active_addr[8] .power_up = "low";

cycloneive_lcell_comb \Selector108~0 (
	.dataa(\m_addr[3]~0_combout ),
	.datab(\active_addr[8]~q ),
	.datac(\WideOr9~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector108~0_combout ),
	.cout());
defparam \Selector108~0 .lut_mask = 16'hDEFF;
defparam \Selector108~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector108~1 (
	.dataa(\active_addr[19]~q ),
	.datab(\m_addr[3]~0_combout ),
	.datac(\Selector108~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[44]~24_combout ),
	.cin(gnd),
	.combout(\Selector108~1_combout ),
	.cout());
defparam \Selector108~1 .lut_mask = 16'hFFBE;
defparam \Selector108~1 .sum_lutc_input = "datac";

dffeas \active_addr[9] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[45]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_addr[9]~q ),
	.prn(vcc));
defparam \active_addr[9] .is_wysiwyg = "true";
defparam \active_addr[9] .power_up = "low";

cycloneive_lcell_comb \Selector107~0 (
	.dataa(\WideOr9~0_combout ),
	.datab(\active_addr[20]~q ),
	.datac(\m_addr[3]~0_combout ),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector107~0_combout ),
	.cout());
defparam \Selector107~0 .lut_mask = 16'hDEFF;
defparam \Selector107~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector107~1 (
	.dataa(\active_addr[9]~q ),
	.datab(\WideOr9~0_combout ),
	.datac(\Selector107~0_combout ),
	.datad(\the_final_project_soc_sdram_input_efifo_module|rd_data[45]~25_combout ),
	.cin(gnd),
	.combout(\Selector107~1_combout ),
	.cout());
defparam \Selector107~1 .lut_mask = 16'hFFBE;
defparam \Selector107~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\pending~combout ),
	.datab(\f_pop~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'h7777;
defparam \always5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector106~2 (
	.dataa(\active_addr[21]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector106~2_combout ),
	.cout());
defparam \Selector106~2 .lut_mask = 16'h88BB;
defparam \Selector106~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector106~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector106~2_combout ),
	.cin(gnd),
	.combout(\Selector106~3_combout ),
	.cout());
defparam \Selector106~3 .lut_mask = 16'hFFF7;
defparam \Selector106~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector105~2 (
	.dataa(\active_addr[22]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector105~2_combout ),
	.cout());
defparam \Selector105~2 .lut_mask = 16'h88BB;
defparam \Selector105~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector105~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector105~2_combout ),
	.cin(gnd),
	.combout(\Selector105~3_combout ),
	.cout());
defparam \Selector105~3 .lut_mask = 16'hFFF7;
defparam \Selector105~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector104~2 (
	.dataa(\active_addr[23]~q ),
	.datab(\m_state.000000010~q ),
	.datac(gnd),
	.datad(\i_addr[12]~q ),
	.cin(gnd),
	.combout(\Selector104~2_combout ),
	.cout());
defparam \Selector104~2 .lut_mask = 16'h88BB;
defparam \Selector104~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector104~3 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.001000000~q ),
	.datad(\Selector104~2_combout ),
	.cin(gnd),
	.combout(\Selector104~3_combout ),
	.cout());
defparam \Selector104~3 .lut_mask = 16'hFFF7;
defparam \Selector104~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector118~0 (
	.dataa(\active_addr[10]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[46]~0_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector118~0_combout ),
	.cout());
defparam \Selector118~0 .lut_mask = 16'hEFFE;
defparam \Selector118~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr16~0 (
	.dataa(\m_state.000001000~q ),
	.datab(\m_state.000010000~q ),
	.datac(\m_state.000000010~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr16~0_combout ),
	.cout());
defparam \WideOr16~0 .lut_mask = 16'hFEFE;
defparam \WideOr16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector117~0 (
	.dataa(\active_addr[24]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[60]~2_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector117~0_combout ),
	.cout());
defparam \Selector117~0 .lut_mask = 16'hEFFE;
defparam \Selector117~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\i_state.001~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[1]~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFFF7;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \i_cmd[1] (
	.clk(wire_pll7_clk_0),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[1]~q ),
	.prn(vcc));
defparam \i_cmd[1] .is_wysiwyg = "true";
defparam \i_cmd[1] .power_up = "low";

cycloneive_lcell_comb \Selector21~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[1]~q ),
	.datac(\m_state.000000001~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
defparam \Selector21~0 .lut_mask = 16'hDFD5;
defparam \Selector21~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector21~1 (
	.dataa(\always5~0_combout ),
	.datab(\WideOr9~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\Selector21~0_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
defparam \Selector21~1 .lut_mask = 16'hFFB8;
defparam \Selector21~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\i_state.101~q ),
	.datab(gnd),
	.datac(\i_cmd[3]~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFFF5;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \i_cmd[3] (
	.clk(wire_pll7_clk_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[3]~q ),
	.prn(vcc));
defparam \i_cmd[3] .is_wysiwyg = "true";
defparam \i_cmd[3] .power_up = "low";

cycloneive_lcell_comb \Selector19~0 (
	.dataa(\init_done~q ),
	.datab(\i_cmd[3]~q ),
	.datac(\refresh_request~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
defparam \Selector19~0 .lut_mask = 16'h27FF;
defparam \Selector19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~1 (
	.dataa(\m_state.000000001~q ),
	.datab(\m_state.001000000~q ),
	.datac(\m_state.000000100~q ),
	.datad(\m_state.010000000~q ),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
defparam \Selector19~1 .lut_mask = 16'hBFFF;
defparam \Selector19~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~2 (
	.dataa(\m_state.001000000~q ),
	.datab(\m_state.000000100~q ),
	.datac(\refresh_request~q ),
	.datad(\m_next.010000000~q ),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
defparam \Selector19~2 .lut_mask = 16'hEFFF;
defparam \Selector19~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~3 (
	.dataa(\Selector19~0_combout ),
	.datab(\active_cs_n~q ),
	.datac(\Selector19~1_combout ),
	.datad(\Selector19~2_combout ),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
defparam \Selector19~3 .lut_mask = 16'h7FFF;
defparam \Selector19~3 .sum_lutc_input = "datac";

dffeas \active_dqm[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[32]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[0]~q ),
	.prn(vcc));
defparam \active_dqm[0] .is_wysiwyg = "true";
defparam \active_dqm[0] .power_up = "low";

cycloneive_lcell_comb \Selector154~0 (
	.dataa(\active_dqm[0]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[32]~26_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector154~0_combout ),
	.cout());
defparam \Selector154~0 .lut_mask = 16'hEFFE;
defparam \Selector154~0 .sum_lutc_input = "datac";

dffeas \active_dqm[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[33]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[1]~q ),
	.prn(vcc));
defparam \active_dqm[1] .is_wysiwyg = "true";
defparam \active_dqm[1] .power_up = "low";

cycloneive_lcell_comb \Selector153~0 (
	.dataa(\active_dqm[1]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[33]~27_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector153~0_combout ),
	.cout());
defparam \Selector153~0 .lut_mask = 16'hEFFE;
defparam \Selector153~0 .sum_lutc_input = "datac";

dffeas \active_dqm[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[34]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[2]~q ),
	.prn(vcc));
defparam \active_dqm[2] .is_wysiwyg = "true";
defparam \active_dqm[2] .power_up = "low";

cycloneive_lcell_comb \Selector152~0 (
	.dataa(\active_dqm[2]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[34]~28_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector152~0_combout ),
	.cout());
defparam \Selector152~0 .lut_mask = 16'hEFFE;
defparam \Selector152~0 .sum_lutc_input = "datac";

dffeas \active_dqm[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[35]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_dqm[3]~q ),
	.prn(vcc));
defparam \active_dqm[3] .is_wysiwyg = "true";
defparam \active_dqm[3] .power_up = "low";

cycloneive_lcell_comb \Selector151~0 (
	.dataa(\active_dqm[3]~q ),
	.datab(\the_final_project_soc_sdram_input_efifo_module|rd_data[35]~29_combout ),
	.datac(\f_select~combout ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector151~0_combout ),
	.cout());
defparam \Selector151~0 .lut_mask = 16'hEFFE;
defparam \Selector151~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\i_state.011~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[2]~q ),
	.datad(\i_state.000~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFFF7;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \i_cmd[2] (
	.clk(wire_pll7_clk_0),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[2]~q ),
	.prn(vcc));
defparam \i_cmd[2] .is_wysiwyg = "true";
defparam \i_cmd[2] .power_up = "low";

cycloneive_lcell_comb \Selector20~0 (
	.dataa(\WideOr8~0_combout ),
	.datab(\init_done~q ),
	.datac(\i_cmd[2]~q ),
	.datad(\m_state.000000001~q ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
defparam \Selector20~0 .lut_mask = 16'hF377;
defparam \Selector20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\i_state.010~q ),
	.datab(\i_state.101~q ),
	.datac(\i_cmd[0]~q ),
	.datad(\WideOr6~0_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFFF7;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \i_cmd[0] (
	.clk(wire_pll7_clk_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_cmd[0]~q ),
	.prn(vcc));
defparam \i_cmd[0] .is_wysiwyg = "true";
defparam \i_cmd[0] .power_up = "low";

cycloneive_lcell_comb \Selector22~0 (
	.dataa(\m_state.000000001~q ),
	.datab(\m_state.001000000~q ),
	.datac(\init_done~q ),
	.datad(\i_cmd[0]~q ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
defparam \Selector22~0 .lut_mask = 16'hDF8F;
defparam \Selector22~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector22~1 (
	.dataa(\m_state.000010000~q ),
	.datab(\always5~0_combout ),
	.datac(\m_state.000000001~q ),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
defparam \Selector22~1 .lut_mask = 16'hFFD8;
defparam \Selector22~1 .sum_lutc_input = "datac";

dffeas \active_data[0] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[0]~q ),
	.prn(vcc));
defparam \active_data[0] .is_wysiwyg = "true";
defparam \active_data[0] .power_up = "low";

cycloneive_lcell_comb \Selector150~0 (
	.dataa(\active_data[0]~q ),
	.datab(m_data_0),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector150~0_combout ),
	.cout());
defparam \Selector150~0 .lut_mask = 16'hEFFE;
defparam \Selector150~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m_data[3]~0 (
	.dataa(\f_pop~q ),
	.datab(\m_state.000010000~q ),
	.datac(gnd),
	.datad(\pending~combout ),
	.cin(gnd),
	.combout(\m_data[3]~0_combout ),
	.cout());
defparam \m_data[3]~0 .lut_mask = 16'hEEFF;
defparam \m_data[3]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector150~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[0]~30_combout ),
	.datab(\Selector150~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector150~1_combout ),
	.cout());
defparam \Selector150~1 .lut_mask = 16'hAACC;
defparam \Selector150~1 .sum_lutc_input = "datac";

dffeas \active_data[1] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[1]~q ),
	.prn(vcc));
defparam \active_data[1] .is_wysiwyg = "true";
defparam \active_data[1] .power_up = "low";

cycloneive_lcell_comb \Selector149~0 (
	.dataa(\active_data[1]~q ),
	.datab(m_data_1),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector149~0_combout ),
	.cout());
defparam \Selector149~0 .lut_mask = 16'hEFFE;
defparam \Selector149~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector149~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[1]~31_combout ),
	.datab(\Selector149~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector149~1_combout ),
	.cout());
defparam \Selector149~1 .lut_mask = 16'hAACC;
defparam \Selector149~1 .sum_lutc_input = "datac";

dffeas \active_data[2] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[2]~q ),
	.prn(vcc));
defparam \active_data[2] .is_wysiwyg = "true";
defparam \active_data[2] .power_up = "low";

cycloneive_lcell_comb \Selector148~0 (
	.dataa(\active_data[2]~q ),
	.datab(m_data_2),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector148~0_combout ),
	.cout());
defparam \Selector148~0 .lut_mask = 16'hEFFE;
defparam \Selector148~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector148~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[2]~32_combout ),
	.datab(\Selector148~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector148~1_combout ),
	.cout());
defparam \Selector148~1 .lut_mask = 16'hAACC;
defparam \Selector148~1 .sum_lutc_input = "datac";

dffeas \active_data[3] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[3]~q ),
	.prn(vcc));
defparam \active_data[3] .is_wysiwyg = "true";
defparam \active_data[3] .power_up = "low";

cycloneive_lcell_comb \Selector147~0 (
	.dataa(\active_data[3]~q ),
	.datab(m_data_3),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector147~0_combout ),
	.cout());
defparam \Selector147~0 .lut_mask = 16'hEFFE;
defparam \Selector147~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector147~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[3]~33_combout ),
	.datab(\Selector147~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector147~1_combout ),
	.cout());
defparam \Selector147~1 .lut_mask = 16'hAACC;
defparam \Selector147~1 .sum_lutc_input = "datac";

dffeas \active_data[4] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[4]~q ),
	.prn(vcc));
defparam \active_data[4] .is_wysiwyg = "true";
defparam \active_data[4] .power_up = "low";

cycloneive_lcell_comb \Selector146~0 (
	.dataa(\active_data[4]~q ),
	.datab(m_data_4),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector146~0_combout ),
	.cout());
defparam \Selector146~0 .lut_mask = 16'hEFFE;
defparam \Selector146~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector146~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[4]~34_combout ),
	.datab(\Selector146~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector146~1_combout ),
	.cout());
defparam \Selector146~1 .lut_mask = 16'hAACC;
defparam \Selector146~1 .sum_lutc_input = "datac";

dffeas \active_data[5] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[5]~q ),
	.prn(vcc));
defparam \active_data[5] .is_wysiwyg = "true";
defparam \active_data[5] .power_up = "low";

cycloneive_lcell_comb \Selector145~0 (
	.dataa(\active_data[5]~q ),
	.datab(m_data_5),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector145~0_combout ),
	.cout());
defparam \Selector145~0 .lut_mask = 16'hEFFE;
defparam \Selector145~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector145~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[5]~35_combout ),
	.datab(\Selector145~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector145~1_combout ),
	.cout());
defparam \Selector145~1 .lut_mask = 16'hAACC;
defparam \Selector145~1 .sum_lutc_input = "datac";

dffeas \active_data[6] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[6]~q ),
	.prn(vcc));
defparam \active_data[6] .is_wysiwyg = "true";
defparam \active_data[6] .power_up = "low";

cycloneive_lcell_comb \Selector144~0 (
	.dataa(\active_data[6]~q ),
	.datab(m_data_6),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector144~0_combout ),
	.cout());
defparam \Selector144~0 .lut_mask = 16'hEFFE;
defparam \Selector144~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector144~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[6]~36_combout ),
	.datab(\Selector144~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector144~1_combout ),
	.cout());
defparam \Selector144~1 .lut_mask = 16'hAACC;
defparam \Selector144~1 .sum_lutc_input = "datac";

dffeas \active_data[7] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[7]~q ),
	.prn(vcc));
defparam \active_data[7] .is_wysiwyg = "true";
defparam \active_data[7] .power_up = "low";

cycloneive_lcell_comb \Selector143~0 (
	.dataa(\active_data[7]~q ),
	.datab(m_data_7),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector143~0_combout ),
	.cout());
defparam \Selector143~0 .lut_mask = 16'hEFFE;
defparam \Selector143~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector143~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[7]~37_combout ),
	.datab(\Selector143~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector143~1_combout ),
	.cout());
defparam \Selector143~1 .lut_mask = 16'hAACC;
defparam \Selector143~1 .sum_lutc_input = "datac";

dffeas \active_data[8] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[8]~q ),
	.prn(vcc));
defparam \active_data[8] .is_wysiwyg = "true";
defparam \active_data[8] .power_up = "low";

cycloneive_lcell_comb \Selector142~0 (
	.dataa(\active_data[8]~q ),
	.datab(m_data_8),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector142~0_combout ),
	.cout());
defparam \Selector142~0 .lut_mask = 16'hEFFE;
defparam \Selector142~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector142~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[8]~38_combout ),
	.datab(\Selector142~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector142~1_combout ),
	.cout());
defparam \Selector142~1 .lut_mask = 16'hAACC;
defparam \Selector142~1 .sum_lutc_input = "datac";

dffeas \active_data[9] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[9]~q ),
	.prn(vcc));
defparam \active_data[9] .is_wysiwyg = "true";
defparam \active_data[9] .power_up = "low";

cycloneive_lcell_comb \Selector141~0 (
	.dataa(\active_data[9]~q ),
	.datab(m_data_9),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector141~0_combout ),
	.cout());
defparam \Selector141~0 .lut_mask = 16'hEFFE;
defparam \Selector141~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector141~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[9]~39_combout ),
	.datab(\Selector141~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector141~1_combout ),
	.cout());
defparam \Selector141~1 .lut_mask = 16'hAACC;
defparam \Selector141~1 .sum_lutc_input = "datac";

dffeas \active_data[10] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[10]~q ),
	.prn(vcc));
defparam \active_data[10] .is_wysiwyg = "true";
defparam \active_data[10] .power_up = "low";

cycloneive_lcell_comb \Selector140~0 (
	.dataa(\active_data[10]~q ),
	.datab(m_data_10),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector140~0_combout ),
	.cout());
defparam \Selector140~0 .lut_mask = 16'hEFFE;
defparam \Selector140~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector140~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[10]~40_combout ),
	.datab(\Selector140~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector140~1_combout ),
	.cout());
defparam \Selector140~1 .lut_mask = 16'hAACC;
defparam \Selector140~1 .sum_lutc_input = "datac";

dffeas \active_data[11] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[11]~q ),
	.prn(vcc));
defparam \active_data[11] .is_wysiwyg = "true";
defparam \active_data[11] .power_up = "low";

cycloneive_lcell_comb \Selector139~0 (
	.dataa(\active_data[11]~q ),
	.datab(m_data_11),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector139~0_combout ),
	.cout());
defparam \Selector139~0 .lut_mask = 16'hEFFE;
defparam \Selector139~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector139~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[11]~41_combout ),
	.datab(\Selector139~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector139~1_combout ),
	.cout());
defparam \Selector139~1 .lut_mask = 16'hAACC;
defparam \Selector139~1 .sum_lutc_input = "datac";

dffeas \active_data[12] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[12]~q ),
	.prn(vcc));
defparam \active_data[12] .is_wysiwyg = "true";
defparam \active_data[12] .power_up = "low";

cycloneive_lcell_comb \Selector138~0 (
	.dataa(\active_data[12]~q ),
	.datab(m_data_12),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector138~0_combout ),
	.cout());
defparam \Selector138~0 .lut_mask = 16'hEFFE;
defparam \Selector138~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector138~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[12]~42_combout ),
	.datab(\Selector138~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector138~1_combout ),
	.cout());
defparam \Selector138~1 .lut_mask = 16'hAACC;
defparam \Selector138~1 .sum_lutc_input = "datac";

dffeas \active_data[13] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[13]~q ),
	.prn(vcc));
defparam \active_data[13] .is_wysiwyg = "true";
defparam \active_data[13] .power_up = "low";

cycloneive_lcell_comb \Selector137~0 (
	.dataa(\active_data[13]~q ),
	.datab(m_data_13),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector137~0_combout ),
	.cout());
defparam \Selector137~0 .lut_mask = 16'hEFFE;
defparam \Selector137~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector137~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[13]~43_combout ),
	.datab(\Selector137~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector137~1_combout ),
	.cout());
defparam \Selector137~1 .lut_mask = 16'hAACC;
defparam \Selector137~1 .sum_lutc_input = "datac";

dffeas \active_data[14] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[14]~q ),
	.prn(vcc));
defparam \active_data[14] .is_wysiwyg = "true";
defparam \active_data[14] .power_up = "low";

cycloneive_lcell_comb \Selector136~0 (
	.dataa(\active_data[14]~q ),
	.datab(m_data_14),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector136~0_combout ),
	.cout());
defparam \Selector136~0 .lut_mask = 16'hEFFE;
defparam \Selector136~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector136~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[14]~44_combout ),
	.datab(\Selector136~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector136~1_combout ),
	.cout());
defparam \Selector136~1 .lut_mask = 16'hAACC;
defparam \Selector136~1 .sum_lutc_input = "datac";

dffeas \active_data[15] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[15]~q ),
	.prn(vcc));
defparam \active_data[15] .is_wysiwyg = "true";
defparam \active_data[15] .power_up = "low";

cycloneive_lcell_comb \Selector135~0 (
	.dataa(\active_data[15]~q ),
	.datab(m_data_15),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector135~0_combout ),
	.cout());
defparam \Selector135~0 .lut_mask = 16'hEFFE;
defparam \Selector135~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector135~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[15]~45_combout ),
	.datab(\Selector135~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector135~1_combout ),
	.cout());
defparam \Selector135~1 .lut_mask = 16'hAACC;
defparam \Selector135~1 .sum_lutc_input = "datac";

dffeas \active_data[16] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[16]~q ),
	.prn(vcc));
defparam \active_data[16] .is_wysiwyg = "true";
defparam \active_data[16] .power_up = "low";

cycloneive_lcell_comb \Selector134~0 (
	.dataa(\active_data[16]~q ),
	.datab(m_data_16),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector134~0_combout ),
	.cout());
defparam \Selector134~0 .lut_mask = 16'hEFFE;
defparam \Selector134~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector134~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[16]~46_combout ),
	.datab(\Selector134~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector134~1_combout ),
	.cout());
defparam \Selector134~1 .lut_mask = 16'hAACC;
defparam \Selector134~1 .sum_lutc_input = "datac";

dffeas \active_data[17] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[17]~q ),
	.prn(vcc));
defparam \active_data[17] .is_wysiwyg = "true";
defparam \active_data[17] .power_up = "low";

cycloneive_lcell_comb \Selector133~0 (
	.dataa(\active_data[17]~q ),
	.datab(m_data_17),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector133~0_combout ),
	.cout());
defparam \Selector133~0 .lut_mask = 16'hEFFE;
defparam \Selector133~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector133~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[17]~47_combout ),
	.datab(\Selector133~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector133~1_combout ),
	.cout());
defparam \Selector133~1 .lut_mask = 16'hAACC;
defparam \Selector133~1 .sum_lutc_input = "datac";

dffeas \active_data[18] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[18]~q ),
	.prn(vcc));
defparam \active_data[18] .is_wysiwyg = "true";
defparam \active_data[18] .power_up = "low";

cycloneive_lcell_comb \Selector132~0 (
	.dataa(\active_data[18]~q ),
	.datab(m_data_18),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector132~0_combout ),
	.cout());
defparam \Selector132~0 .lut_mask = 16'hEFFE;
defparam \Selector132~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector132~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[18]~48_combout ),
	.datab(\Selector132~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector132~1_combout ),
	.cout());
defparam \Selector132~1 .lut_mask = 16'hAACC;
defparam \Selector132~1 .sum_lutc_input = "datac";

dffeas \active_data[19] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[19]~q ),
	.prn(vcc));
defparam \active_data[19] .is_wysiwyg = "true";
defparam \active_data[19] .power_up = "low";

cycloneive_lcell_comb \Selector131~0 (
	.dataa(\active_data[19]~q ),
	.datab(m_data_19),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector131~0_combout ),
	.cout());
defparam \Selector131~0 .lut_mask = 16'hEFFE;
defparam \Selector131~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector131~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[19]~49_combout ),
	.datab(\Selector131~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector131~1_combout ),
	.cout());
defparam \Selector131~1 .lut_mask = 16'hAACC;
defparam \Selector131~1 .sum_lutc_input = "datac";

dffeas \active_data[20] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[20]~q ),
	.prn(vcc));
defparam \active_data[20] .is_wysiwyg = "true";
defparam \active_data[20] .power_up = "low";

cycloneive_lcell_comb \Selector130~0 (
	.dataa(\active_data[20]~q ),
	.datab(m_data_20),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector130~0_combout ),
	.cout());
defparam \Selector130~0 .lut_mask = 16'hEFFE;
defparam \Selector130~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector130~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[20]~50_combout ),
	.datab(\Selector130~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector130~1_combout ),
	.cout());
defparam \Selector130~1 .lut_mask = 16'hAACC;
defparam \Selector130~1 .sum_lutc_input = "datac";

dffeas \active_data[21] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[21]~q ),
	.prn(vcc));
defparam \active_data[21] .is_wysiwyg = "true";
defparam \active_data[21] .power_up = "low";

cycloneive_lcell_comb \Selector129~0 (
	.dataa(\active_data[21]~q ),
	.datab(m_data_21),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector129~0_combout ),
	.cout());
defparam \Selector129~0 .lut_mask = 16'hEFFE;
defparam \Selector129~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector129~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[21]~51_combout ),
	.datab(\Selector129~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector129~1_combout ),
	.cout());
defparam \Selector129~1 .lut_mask = 16'hAACC;
defparam \Selector129~1 .sum_lutc_input = "datac";

dffeas \active_data[22] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[22]~q ),
	.prn(vcc));
defparam \active_data[22] .is_wysiwyg = "true";
defparam \active_data[22] .power_up = "low";

cycloneive_lcell_comb \Selector128~0 (
	.dataa(\active_data[22]~q ),
	.datab(m_data_22),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector128~0_combout ),
	.cout());
defparam \Selector128~0 .lut_mask = 16'hEFFE;
defparam \Selector128~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector128~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[22]~52_combout ),
	.datab(\Selector128~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector128~1_combout ),
	.cout());
defparam \Selector128~1 .lut_mask = 16'hAACC;
defparam \Selector128~1 .sum_lutc_input = "datac";

dffeas \active_data[23] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[23]~q ),
	.prn(vcc));
defparam \active_data[23] .is_wysiwyg = "true";
defparam \active_data[23] .power_up = "low";

cycloneive_lcell_comb \Selector127~0 (
	.dataa(\active_data[23]~q ),
	.datab(m_data_23),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector127~0_combout ),
	.cout());
defparam \Selector127~0 .lut_mask = 16'hEFFE;
defparam \Selector127~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector127~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[23]~53_combout ),
	.datab(\Selector127~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector127~1_combout ),
	.cout());
defparam \Selector127~1 .lut_mask = 16'hAACC;
defparam \Selector127~1 .sum_lutc_input = "datac";

dffeas \active_data[24] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[24]~q ),
	.prn(vcc));
defparam \active_data[24] .is_wysiwyg = "true";
defparam \active_data[24] .power_up = "low";

cycloneive_lcell_comb \Selector126~0 (
	.dataa(\active_data[24]~q ),
	.datab(m_data_24),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector126~0_combout ),
	.cout());
defparam \Selector126~0 .lut_mask = 16'hEFFE;
defparam \Selector126~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector126~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[24]~54_combout ),
	.datab(\Selector126~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector126~1_combout ),
	.cout());
defparam \Selector126~1 .lut_mask = 16'hAACC;
defparam \Selector126~1 .sum_lutc_input = "datac";

dffeas \active_data[25] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[25]~q ),
	.prn(vcc));
defparam \active_data[25] .is_wysiwyg = "true";
defparam \active_data[25] .power_up = "low";

cycloneive_lcell_comb \Selector125~0 (
	.dataa(\active_data[25]~q ),
	.datab(m_data_25),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector125~0_combout ),
	.cout());
defparam \Selector125~0 .lut_mask = 16'hEFFE;
defparam \Selector125~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector125~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[25]~55_combout ),
	.datab(\Selector125~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector125~1_combout ),
	.cout());
defparam \Selector125~1 .lut_mask = 16'hAACC;
defparam \Selector125~1 .sum_lutc_input = "datac";

dffeas \active_data[26] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[26]~q ),
	.prn(vcc));
defparam \active_data[26] .is_wysiwyg = "true";
defparam \active_data[26] .power_up = "low";

cycloneive_lcell_comb \Selector124~0 (
	.dataa(\active_data[26]~q ),
	.datab(m_data_26),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector124~0_combout ),
	.cout());
defparam \Selector124~0 .lut_mask = 16'hEFFE;
defparam \Selector124~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector124~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[26]~56_combout ),
	.datab(\Selector124~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector124~1_combout ),
	.cout());
defparam \Selector124~1 .lut_mask = 16'hAACC;
defparam \Selector124~1 .sum_lutc_input = "datac";

dffeas \active_data[27] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[27]~q ),
	.prn(vcc));
defparam \active_data[27] .is_wysiwyg = "true";
defparam \active_data[27] .power_up = "low";

cycloneive_lcell_comb \Selector123~0 (
	.dataa(\active_data[27]~q ),
	.datab(m_data_27),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector123~0_combout ),
	.cout());
defparam \Selector123~0 .lut_mask = 16'hEFFE;
defparam \Selector123~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector123~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[27]~57_combout ),
	.datab(\Selector123~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector123~1_combout ),
	.cout());
defparam \Selector123~1 .lut_mask = 16'hAACC;
defparam \Selector123~1 .sum_lutc_input = "datac";

dffeas \active_data[28] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[28]~q ),
	.prn(vcc));
defparam \active_data[28] .is_wysiwyg = "true";
defparam \active_data[28] .power_up = "low";

cycloneive_lcell_comb \Selector122~0 (
	.dataa(\active_data[28]~q ),
	.datab(m_data_28),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector122~0_combout ),
	.cout());
defparam \Selector122~0 .lut_mask = 16'hEFFE;
defparam \Selector122~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector122~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[28]~58_combout ),
	.datab(\Selector122~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector122~1_combout ),
	.cout());
defparam \Selector122~1 .lut_mask = 16'hAACC;
defparam \Selector122~1 .sum_lutc_input = "datac";

dffeas \active_data[29] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[29]~q ),
	.prn(vcc));
defparam \active_data[29] .is_wysiwyg = "true";
defparam \active_data[29] .power_up = "low";

cycloneive_lcell_comb \Selector121~0 (
	.dataa(\active_data[29]~q ),
	.datab(m_data_29),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector121~0_combout ),
	.cout());
defparam \Selector121~0 .lut_mask = 16'hEFFE;
defparam \Selector121~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector121~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[29]~59_combout ),
	.datab(\Selector121~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector121~1_combout ),
	.cout());
defparam \Selector121~1 .lut_mask = 16'hAACC;
defparam \Selector121~1 .sum_lutc_input = "datac";

dffeas \active_data[30] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[30]~q ),
	.prn(vcc));
defparam \active_data[30] .is_wysiwyg = "true";
defparam \active_data[30] .power_up = "low";

cycloneive_lcell_comb \Selector120~0 (
	.dataa(\active_data[30]~q ),
	.datab(m_data_30),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector120~0_combout ),
	.cout());
defparam \Selector120~0 .lut_mask = 16'hEFFE;
defparam \Selector120~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector120~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[30]~60_combout ),
	.datab(\Selector120~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector120~1_combout ),
	.cout());
defparam \Selector120~1 .lut_mask = 16'hAACC;
defparam \Selector120~1 .sum_lutc_input = "datac";

dffeas \active_data[31] (
	.clk(wire_pll7_clk_0),
	.d(\the_final_project_soc_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\active_rnw~3_combout ),
	.q(\active_data[31]~q ),
	.prn(vcc));
defparam \active_data[31] .is_wysiwyg = "true";
defparam \active_data[31] .power_up = "low";

cycloneive_lcell_comb \Selector119~0 (
	.dataa(\active_data[31]~q ),
	.datab(m_data_31),
	.datac(\m_state.000010000~q ),
	.datad(\m_state.000000010~q ),
	.cin(gnd),
	.combout(\Selector119~0_combout ),
	.cout());
defparam \Selector119~0 .lut_mask = 16'hEFFE;
defparam \Selector119~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector119~1 (
	.dataa(\the_final_project_soc_sdram_input_efifo_module|rd_data[31]~61_combout ),
	.datab(\Selector119~0_combout ),
	.datac(gnd),
	.datad(\m_data[3]~0_combout ),
	.cin(gnd),
	.combout(\Selector119~1_combout ),
	.cout());
defparam \Selector119~1 .lut_mask = 16'hAACC;
defparam \Selector119~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~0 (
	.dataa(m_cmd_1),
	.datab(gnd),
	.datac(m_cmd_2),
	.datad(m_cmd_0),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hAFFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

dffeas \rd_valid[0] (
	.clk(wire_pll7_clk_0),
	.d(\Equal4~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[0]~q ),
	.prn(vcc));
defparam \rd_valid[0] .is_wysiwyg = "true";
defparam \rd_valid[0] .power_up = "low";

dffeas \rd_valid[1] (
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[1]~q ),
	.prn(vcc));
defparam \rd_valid[1] .is_wysiwyg = "true";
defparam \rd_valid[1] .power_up = "low";

dffeas \rd_valid[2] (
	.clk(wire_pll7_clk_0),
	.d(\rd_valid[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_valid[2]~q ),
	.prn(vcc));
defparam \rd_valid[2] .is_wysiwyg = "true";
defparam \rd_valid[2] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_sdram_input_efifo_module (
	clk,
	f_pop,
	entries_1,
	entries_0,
	Equal1,
	rd_data_46,
	rd_data_61,
	rd_data_60,
	rd_data_47,
	rd_data_49,
	rd_data_48,
	rd_data_51,
	rd_data_50,
	rd_data_53,
	rd_data_52,
	rd_data_55,
	rd_data_54,
	rd_data_57,
	rd_data_56,
	rd_data_59,
	rd_data_58,
	pending,
	rd_data_36,
	reset_n,
	rd_data_37,
	rd_data_38,
	rd_data_39,
	rd_data_40,
	rd_data_41,
	f_select,
	rd_data_42,
	rd_data_43,
	rd_data_44,
	rd_data_45,
	rd_data_32,
	rd_data_33,
	rd_data_34,
	rd_data_35,
	last_cycle,
	WideOr1,
	src_payload,
	src_data_68,
	src_data_48,
	src_data_62,
	src_data_49,
	src_data_51,
	src_data_50,
	src_data_53,
	src_data_52,
	src_data_55,
	src_data_54,
	src_data_57,
	src_data_56,
	src_data_59,
	src_data_58,
	src_data_61,
	src_data_60,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	comb,
	comb1,
	comb2,
	comb3,
	rd_data_0,
	rd_data_1,
	rd_data_2,
	rd_data_3,
	rd_data_4,
	rd_data_5,
	rd_data_6,
	rd_data_7,
	rd_data_8,
	rd_data_9,
	rd_data_10,
	rd_data_11,
	rd_data_12,
	rd_data_13,
	rd_data_14,
	rd_data_15,
	rd_data_16,
	rd_data_17,
	rd_data_18,
	rd_data_19,
	rd_data_20,
	rd_data_21,
	rd_data_22,
	rd_data_23,
	rd_data_24,
	rd_data_25,
	rd_data_26,
	rd_data_27,
	rd_data_28,
	rd_data_29,
	rd_data_30,
	rd_data_31,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	f_pop;
output 	entries_1;
output 	entries_0;
output 	Equal1;
output 	rd_data_46;
output 	rd_data_61;
output 	rd_data_60;
output 	rd_data_47;
output 	rd_data_49;
output 	rd_data_48;
output 	rd_data_51;
output 	rd_data_50;
output 	rd_data_53;
output 	rd_data_52;
output 	rd_data_55;
output 	rd_data_54;
output 	rd_data_57;
output 	rd_data_56;
output 	rd_data_59;
output 	rd_data_58;
input 	pending;
output 	rd_data_36;
input 	reset_n;
output 	rd_data_37;
output 	rd_data_38;
output 	rd_data_39;
output 	rd_data_40;
output 	rd_data_41;
input 	f_select;
output 	rd_data_42;
output 	rd_data_43;
output 	rd_data_44;
output 	rd_data_45;
output 	rd_data_32;
output 	rd_data_33;
output 	rd_data_34;
output 	rd_data_35;
input 	last_cycle;
input 	WideOr1;
input 	src_payload;
input 	src_data_68;
input 	src_data_48;
input 	src_data_62;
input 	src_data_49;
input 	src_data_51;
input 	src_data_50;
input 	src_data_53;
input 	src_data_52;
input 	src_data_55;
input 	src_data_54;
input 	src_data_57;
input 	src_data_56;
input 	src_data_59;
input 	src_data_58;
input 	src_data_61;
input 	src_data_60;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	comb;
input 	comb1;
input 	comb2;
input 	comb3;
output 	rd_data_0;
output 	rd_data_1;
output 	rd_data_2;
output 	rd_data_3;
output 	rd_data_4;
output 	rd_data_5;
output 	rd_data_6;
output 	rd_data_7;
output 	rd_data_8;
output 	rd_data_9;
output 	rd_data_10;
output 	rd_data_11;
output 	rd_data_12;
output 	rd_data_13;
output 	rd_data_14;
output 	rd_data_15;
output 	rd_data_16;
output 	rd_data_17;
output 	rd_data_18;
output 	rd_data_19;
output 	rd_data_20;
output 	rd_data_21;
output 	rd_data_22;
output 	rd_data_23;
output 	rd_data_24;
output 	rd_data_25;
output 	rd_data_26;
output 	rd_data_27;
output 	rd_data_28;
output 	rd_data_29;
output 	rd_data_30;
output 	rd_data_31;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always2~0_combout ;
wire \entries[1]~0_combout ;
wire \entries[0]~1_combout ;
wire \wr_address~0_combout ;
wire \wr_address~q ;
wire \entry_1[61]~0_combout ;
wire \entry_1[46]~q ;
wire \entry_0[61]~0_combout ;
wire \entry_0[46]~q ;
wire \rd_address~0_combout ;
wire \rd_address~q ;
wire \entry_1[61]~q ;
wire \entry_0[61]~q ;
wire \entry_1[60]~q ;
wire \entry_0[60]~q ;
wire \entry_1[47]~q ;
wire \entry_0[47]~q ;
wire \entry_1[49]~q ;
wire \entry_0[49]~q ;
wire \entry_1[48]~q ;
wire \entry_0[48]~q ;
wire \entry_1[51]~q ;
wire \entry_0[51]~q ;
wire \entry_1[50]~q ;
wire \entry_0[50]~q ;
wire \entry_1[53]~q ;
wire \entry_0[53]~q ;
wire \entry_1[52]~q ;
wire \entry_0[52]~q ;
wire \entry_1[55]~q ;
wire \entry_0[55]~q ;
wire \entry_1[54]~q ;
wire \entry_0[54]~q ;
wire \entry_1[57]~q ;
wire \entry_0[57]~q ;
wire \entry_1[56]~q ;
wire \entry_0[56]~q ;
wire \entry_1[59]~q ;
wire \entry_0[59]~q ;
wire \entry_1[58]~q ;
wire \entry_0[58]~q ;
wire \entry_1[36]~q ;
wire \entry_0[36]~q ;
wire \entry_1[37]~q ;
wire \entry_0[37]~q ;
wire \entry_1[38]~q ;
wire \entry_0[38]~q ;
wire \entry_1[39]~q ;
wire \entry_0[39]~q ;
wire \entry_1[40]~q ;
wire \entry_0[40]~q ;
wire \entry_1[41]~q ;
wire \entry_0[41]~q ;
wire \entry_1[42]~q ;
wire \entry_0[42]~q ;
wire \entry_1[43]~q ;
wire \entry_0[43]~q ;
wire \entry_1[44]~q ;
wire \entry_0[44]~q ;
wire \entry_1[45]~q ;
wire \entry_0[45]~q ;
wire \entry_1[32]~q ;
wire \entry_0[32]~q ;
wire \entry_1[33]~q ;
wire \entry_0[33]~q ;
wire \entry_1[34]~q ;
wire \entry_0[34]~q ;
wire \entry_1[35]~q ;
wire \entry_0[35]~q ;
wire \entry_1[0]~q ;
wire \entry_0[0]~q ;
wire \entry_1[1]~q ;
wire \entry_0[1]~q ;
wire \entry_1[2]~q ;
wire \entry_0[2]~q ;
wire \entry_1[3]~q ;
wire \entry_0[3]~q ;
wire \entry_1[4]~q ;
wire \entry_0[4]~q ;
wire \entry_1[5]~q ;
wire \entry_0[5]~q ;
wire \entry_1[6]~q ;
wire \entry_0[6]~q ;
wire \entry_1[7]~q ;
wire \entry_0[7]~q ;
wire \entry_1[8]~q ;
wire \entry_0[8]~q ;
wire \entry_1[9]~q ;
wire \entry_0[9]~q ;
wire \entry_1[10]~q ;
wire \entry_0[10]~q ;
wire \entry_1[11]~q ;
wire \entry_0[11]~q ;
wire \entry_1[12]~q ;
wire \entry_0[12]~q ;
wire \entry_1[13]~q ;
wire \entry_0[13]~q ;
wire \entry_1[14]~q ;
wire \entry_0[14]~q ;
wire \entry_1[15]~q ;
wire \entry_0[15]~q ;
wire \entry_1[16]~q ;
wire \entry_0[16]~q ;
wire \entry_1[17]~q ;
wire \entry_0[17]~q ;
wire \entry_1[18]~q ;
wire \entry_0[18]~q ;
wire \entry_1[19]~q ;
wire \entry_0[19]~q ;
wire \entry_1[20]~q ;
wire \entry_0[20]~q ;
wire \entry_1[21]~q ;
wire \entry_0[21]~q ;
wire \entry_1[22]~q ;
wire \entry_0[22]~q ;
wire \entry_1[23]~q ;
wire \entry_0[23]~q ;
wire \entry_1[24]~q ;
wire \entry_0[24]~q ;
wire \entry_1[25]~q ;
wire \entry_0[25]~q ;
wire \entry_1[26]~q ;
wire \entry_0[26]~q ;
wire \entry_1[27]~q ;
wire \entry_0[27]~q ;
wire \entry_1[28]~q ;
wire \entry_0[28]~q ;
wire \entry_1[29]~q ;
wire \entry_0[29]~q ;
wire \entry_1[30]~q ;
wire \entry_0[30]~q ;
wire \entry_1[31]~q ;
wire \entry_0[31]~q ;


dffeas \entries[1] (
	.clk(clk),
	.d(\entries[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_1),
	.prn(vcc));
defparam \entries[1] .is_wysiwyg = "true";
defparam \entries[1] .power_up = "low";

dffeas \entries[0] (
	.clk(clk),
	.d(\entries[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(entries_0),
	.prn(vcc));
defparam \entries[0] .is_wysiwyg = "true";
defparam \entries[0] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(entries_1),
	.datab(entries_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEEEE;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[46]~0 (
	.dataa(\entry_1[46]~q ),
	.datab(\entry_0[46]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_46),
	.cout());
defparam \rd_data[46]~0 .lut_mask = 16'hAACC;
defparam \rd_data[46]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[61]~1 (
	.dataa(\entry_1[61]~q ),
	.datab(\entry_0[61]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_61),
	.cout());
defparam \rd_data[61]~1 .lut_mask = 16'hAACC;
defparam \rd_data[61]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[60]~2 (
	.dataa(\entry_1[60]~q ),
	.datab(\entry_0[60]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_60),
	.cout());
defparam \rd_data[60]~2 .lut_mask = 16'hAACC;
defparam \rd_data[60]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[47]~3 (
	.dataa(\entry_1[47]~q ),
	.datab(\entry_0[47]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_47),
	.cout());
defparam \rd_data[47]~3 .lut_mask = 16'hAACC;
defparam \rd_data[47]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[49]~4 (
	.dataa(\entry_1[49]~q ),
	.datab(\entry_0[49]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_49),
	.cout());
defparam \rd_data[49]~4 .lut_mask = 16'hAACC;
defparam \rd_data[49]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[48]~5 (
	.dataa(\entry_1[48]~q ),
	.datab(\entry_0[48]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_48),
	.cout());
defparam \rd_data[48]~5 .lut_mask = 16'hAACC;
defparam \rd_data[48]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[51]~6 (
	.dataa(\entry_1[51]~q ),
	.datab(\entry_0[51]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_51),
	.cout());
defparam \rd_data[51]~6 .lut_mask = 16'hAACC;
defparam \rd_data[51]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[50]~7 (
	.dataa(\entry_1[50]~q ),
	.datab(\entry_0[50]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_50),
	.cout());
defparam \rd_data[50]~7 .lut_mask = 16'hAACC;
defparam \rd_data[50]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[53]~8 (
	.dataa(\entry_1[53]~q ),
	.datab(\entry_0[53]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_53),
	.cout());
defparam \rd_data[53]~8 .lut_mask = 16'hAACC;
defparam \rd_data[53]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[52]~9 (
	.dataa(\entry_1[52]~q ),
	.datab(\entry_0[52]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_52),
	.cout());
defparam \rd_data[52]~9 .lut_mask = 16'hAACC;
defparam \rd_data[52]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[55]~10 (
	.dataa(\entry_1[55]~q ),
	.datab(\entry_0[55]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_55),
	.cout());
defparam \rd_data[55]~10 .lut_mask = 16'hAACC;
defparam \rd_data[55]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[54]~11 (
	.dataa(\entry_1[54]~q ),
	.datab(\entry_0[54]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_54),
	.cout());
defparam \rd_data[54]~11 .lut_mask = 16'hAACC;
defparam \rd_data[54]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[57]~12 (
	.dataa(\entry_1[57]~q ),
	.datab(\entry_0[57]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_57),
	.cout());
defparam \rd_data[57]~12 .lut_mask = 16'hAACC;
defparam \rd_data[57]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[56]~13 (
	.dataa(\entry_1[56]~q ),
	.datab(\entry_0[56]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_56),
	.cout());
defparam \rd_data[56]~13 .lut_mask = 16'hAACC;
defparam \rd_data[56]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[59]~14 (
	.dataa(\entry_1[59]~q ),
	.datab(\entry_0[59]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_59),
	.cout());
defparam \rd_data[59]~14 .lut_mask = 16'hAACC;
defparam \rd_data[59]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[58]~15 (
	.dataa(\entry_1[58]~q ),
	.datab(\entry_0[58]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_58),
	.cout());
defparam \rd_data[58]~15 .lut_mask = 16'hAACC;
defparam \rd_data[58]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[36]~16 (
	.dataa(\entry_1[36]~q ),
	.datab(\entry_0[36]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_36),
	.cout());
defparam \rd_data[36]~16 .lut_mask = 16'hAACC;
defparam \rd_data[36]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[37]~17 (
	.dataa(\entry_1[37]~q ),
	.datab(\entry_0[37]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_37),
	.cout());
defparam \rd_data[37]~17 .lut_mask = 16'hAACC;
defparam \rd_data[37]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[38]~18 (
	.dataa(\entry_1[38]~q ),
	.datab(\entry_0[38]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_38),
	.cout());
defparam \rd_data[38]~18 .lut_mask = 16'hAACC;
defparam \rd_data[38]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[39]~19 (
	.dataa(\entry_1[39]~q ),
	.datab(\entry_0[39]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_39),
	.cout());
defparam \rd_data[39]~19 .lut_mask = 16'hAACC;
defparam \rd_data[39]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[40]~20 (
	.dataa(\entry_1[40]~q ),
	.datab(\entry_0[40]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_40),
	.cout());
defparam \rd_data[40]~20 .lut_mask = 16'hAACC;
defparam \rd_data[40]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[41]~21 (
	.dataa(\entry_1[41]~q ),
	.datab(\entry_0[41]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_41),
	.cout());
defparam \rd_data[41]~21 .lut_mask = 16'hAACC;
defparam \rd_data[41]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[42]~22 (
	.dataa(\entry_1[42]~q ),
	.datab(\entry_0[42]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_42),
	.cout());
defparam \rd_data[42]~22 .lut_mask = 16'hAACC;
defparam \rd_data[42]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[43]~23 (
	.dataa(\entry_1[43]~q ),
	.datab(\entry_0[43]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_43),
	.cout());
defparam \rd_data[43]~23 .lut_mask = 16'hAACC;
defparam \rd_data[43]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[44]~24 (
	.dataa(\entry_1[44]~q ),
	.datab(\entry_0[44]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_44),
	.cout());
defparam \rd_data[44]~24 .lut_mask = 16'hAACC;
defparam \rd_data[44]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[45]~25 (
	.dataa(\entry_1[45]~q ),
	.datab(\entry_0[45]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_45),
	.cout());
defparam \rd_data[45]~25 .lut_mask = 16'hAACC;
defparam \rd_data[45]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[32]~26 (
	.dataa(\entry_1[32]~q ),
	.datab(\entry_0[32]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_32),
	.cout());
defparam \rd_data[32]~26 .lut_mask = 16'hAACC;
defparam \rd_data[32]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[33]~27 (
	.dataa(\entry_1[33]~q ),
	.datab(\entry_0[33]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_33),
	.cout());
defparam \rd_data[33]~27 .lut_mask = 16'hAACC;
defparam \rd_data[33]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[34]~28 (
	.dataa(\entry_1[34]~q ),
	.datab(\entry_0[34]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_34),
	.cout());
defparam \rd_data[34]~28 .lut_mask = 16'hAACC;
defparam \rd_data[34]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[35]~29 (
	.dataa(\entry_1[35]~q ),
	.datab(\entry_0[35]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_35),
	.cout());
defparam \rd_data[35]~29 .lut_mask = 16'hAACC;
defparam \rd_data[35]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[0]~30 (
	.dataa(\entry_1[0]~q ),
	.datab(\entry_0[0]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_0),
	.cout());
defparam \rd_data[0]~30 .lut_mask = 16'hAACC;
defparam \rd_data[0]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[1]~31 (
	.dataa(\entry_1[1]~q ),
	.datab(\entry_0[1]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_1),
	.cout());
defparam \rd_data[1]~31 .lut_mask = 16'hAACC;
defparam \rd_data[1]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[2]~32 (
	.dataa(\entry_1[2]~q ),
	.datab(\entry_0[2]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_2),
	.cout());
defparam \rd_data[2]~32 .lut_mask = 16'hAACC;
defparam \rd_data[2]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[3]~33 (
	.dataa(\entry_1[3]~q ),
	.datab(\entry_0[3]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_3),
	.cout());
defparam \rd_data[3]~33 .lut_mask = 16'hAACC;
defparam \rd_data[3]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[4]~34 (
	.dataa(\entry_1[4]~q ),
	.datab(\entry_0[4]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_4),
	.cout());
defparam \rd_data[4]~34 .lut_mask = 16'hAACC;
defparam \rd_data[4]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[5]~35 (
	.dataa(\entry_1[5]~q ),
	.datab(\entry_0[5]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_5),
	.cout());
defparam \rd_data[5]~35 .lut_mask = 16'hAACC;
defparam \rd_data[5]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[6]~36 (
	.dataa(\entry_1[6]~q ),
	.datab(\entry_0[6]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_6),
	.cout());
defparam \rd_data[6]~36 .lut_mask = 16'hAACC;
defparam \rd_data[6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[7]~37 (
	.dataa(\entry_1[7]~q ),
	.datab(\entry_0[7]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_7),
	.cout());
defparam \rd_data[7]~37 .lut_mask = 16'hAACC;
defparam \rd_data[7]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[8]~38 (
	.dataa(\entry_1[8]~q ),
	.datab(\entry_0[8]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_8),
	.cout());
defparam \rd_data[8]~38 .lut_mask = 16'hAACC;
defparam \rd_data[8]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[9]~39 (
	.dataa(\entry_1[9]~q ),
	.datab(\entry_0[9]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_9),
	.cout());
defparam \rd_data[9]~39 .lut_mask = 16'hAACC;
defparam \rd_data[9]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[10]~40 (
	.dataa(\entry_1[10]~q ),
	.datab(\entry_0[10]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_10),
	.cout());
defparam \rd_data[10]~40 .lut_mask = 16'hAACC;
defparam \rd_data[10]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[11]~41 (
	.dataa(\entry_1[11]~q ),
	.datab(\entry_0[11]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_11),
	.cout());
defparam \rd_data[11]~41 .lut_mask = 16'hAACC;
defparam \rd_data[11]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[12]~42 (
	.dataa(\entry_1[12]~q ),
	.datab(\entry_0[12]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_12),
	.cout());
defparam \rd_data[12]~42 .lut_mask = 16'hAACC;
defparam \rd_data[12]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[13]~43 (
	.dataa(\entry_1[13]~q ),
	.datab(\entry_0[13]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_13),
	.cout());
defparam \rd_data[13]~43 .lut_mask = 16'hAACC;
defparam \rd_data[13]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[14]~44 (
	.dataa(\entry_1[14]~q ),
	.datab(\entry_0[14]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_14),
	.cout());
defparam \rd_data[14]~44 .lut_mask = 16'hAACC;
defparam \rd_data[14]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[15]~45 (
	.dataa(\entry_1[15]~q ),
	.datab(\entry_0[15]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_15),
	.cout());
defparam \rd_data[15]~45 .lut_mask = 16'hAACC;
defparam \rd_data[15]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[16]~46 (
	.dataa(\entry_1[16]~q ),
	.datab(\entry_0[16]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_16),
	.cout());
defparam \rd_data[16]~46 .lut_mask = 16'hAACC;
defparam \rd_data[16]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[17]~47 (
	.dataa(\entry_1[17]~q ),
	.datab(\entry_0[17]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_17),
	.cout());
defparam \rd_data[17]~47 .lut_mask = 16'hAACC;
defparam \rd_data[17]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[18]~48 (
	.dataa(\entry_1[18]~q ),
	.datab(\entry_0[18]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_18),
	.cout());
defparam \rd_data[18]~48 .lut_mask = 16'hAACC;
defparam \rd_data[18]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[19]~49 (
	.dataa(\entry_1[19]~q ),
	.datab(\entry_0[19]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_19),
	.cout());
defparam \rd_data[19]~49 .lut_mask = 16'hAACC;
defparam \rd_data[19]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[20]~50 (
	.dataa(\entry_1[20]~q ),
	.datab(\entry_0[20]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_20),
	.cout());
defparam \rd_data[20]~50 .lut_mask = 16'hAACC;
defparam \rd_data[20]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[21]~51 (
	.dataa(\entry_1[21]~q ),
	.datab(\entry_0[21]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_21),
	.cout());
defparam \rd_data[21]~51 .lut_mask = 16'hAACC;
defparam \rd_data[21]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[22]~52 (
	.dataa(\entry_1[22]~q ),
	.datab(\entry_0[22]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_22),
	.cout());
defparam \rd_data[22]~52 .lut_mask = 16'hAACC;
defparam \rd_data[22]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[23]~53 (
	.dataa(\entry_1[23]~q ),
	.datab(\entry_0[23]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_23),
	.cout());
defparam \rd_data[23]~53 .lut_mask = 16'hAACC;
defparam \rd_data[23]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[24]~54 (
	.dataa(\entry_1[24]~q ),
	.datab(\entry_0[24]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_24),
	.cout());
defparam \rd_data[24]~54 .lut_mask = 16'hAACC;
defparam \rd_data[24]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[25]~55 (
	.dataa(\entry_1[25]~q ),
	.datab(\entry_0[25]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_25),
	.cout());
defparam \rd_data[25]~55 .lut_mask = 16'hAACC;
defparam \rd_data[25]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[26]~56 (
	.dataa(\entry_1[26]~q ),
	.datab(\entry_0[26]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_26),
	.cout());
defparam \rd_data[26]~56 .lut_mask = 16'hAACC;
defparam \rd_data[26]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[27]~57 (
	.dataa(\entry_1[27]~q ),
	.datab(\entry_0[27]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_27),
	.cout());
defparam \rd_data[27]~57 .lut_mask = 16'hAACC;
defparam \rd_data[27]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[28]~58 (
	.dataa(\entry_1[28]~q ),
	.datab(\entry_0[28]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_28),
	.cout());
defparam \rd_data[28]~58 .lut_mask = 16'hAACC;
defparam \rd_data[28]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[29]~59 (
	.dataa(\entry_1[29]~q ),
	.datab(\entry_0[29]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_29),
	.cout());
defparam \rd_data[29]~59 .lut_mask = 16'hAACC;
defparam \rd_data[29]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[30]~60 (
	.dataa(\entry_1[30]~q ),
	.datab(\entry_0[30]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_30),
	.cout());
defparam \rd_data[30]~60 .lut_mask = 16'hAACC;
defparam \rd_data[30]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_data[31]~61 (
	.dataa(\entry_1[31]~q ),
	.datab(\entry_0[31]~q ),
	.datac(gnd),
	.datad(\rd_address~q ),
	.cin(gnd),
	.combout(rd_data_31),
	.cout());
defparam \rd_data[31]~61 .lut_mask = 16'hAACC;
defparam \rd_data[31]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(last_cycle),
	.datab(WideOr1),
	.datac(src_payload),
	.datad(src_data_68),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hFFFE;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entries[1]~0 (
	.dataa(entries_1),
	.datab(f_select),
	.datac(entries_0),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\entries[1]~0_combout ),
	.cout());
defparam \entries[1]~0 .lut_mask = 16'h6996;
defparam \entries[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \entries[0]~1 (
	.dataa(f_pop),
	.datab(pending),
	.datac(entries_0),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\entries[0]~1_combout ),
	.cout());
defparam \entries[0]~1 .lut_mask = 16'h6996;
defparam \entries[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_address~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\always2~0_combout ),
	.datad(\wr_address~q ),
	.cin(gnd),
	.combout(\wr_address~0_combout ),
	.cout());
defparam \wr_address~0 .lut_mask = 16'h0FF0;
defparam \wr_address~0 .sum_lutc_input = "datac";

dffeas wr_address(
	.clk(clk),
	.d(\wr_address~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_address~q ),
	.prn(vcc));
defparam wr_address.is_wysiwyg = "true";
defparam wr_address.power_up = "low";

cycloneive_lcell_comb \entry_1[61]~0 (
	.dataa(\always2~0_combout ),
	.datab(\wr_address~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\entry_1[61]~0_combout ),
	.cout());
defparam \entry_1[61]~0 .lut_mask = 16'hEEEE;
defparam \entry_1[61]~0 .sum_lutc_input = "datac";

dffeas \entry_1[46] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[46]~q ),
	.prn(vcc));
defparam \entry_1[46] .is_wysiwyg = "true";
defparam \entry_1[46] .power_up = "low";

cycloneive_lcell_comb \entry_0[61]~0 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wr_address~q ),
	.cin(gnd),
	.combout(\entry_0[61]~0_combout ),
	.cout());
defparam \entry_0[61]~0 .lut_mask = 16'hAAFF;
defparam \entry_0[61]~0 .sum_lutc_input = "datac";

dffeas \entry_0[46] (
	.clk(clk),
	.d(src_data_48),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[46]~q ),
	.prn(vcc));
defparam \entry_0[46] .is_wysiwyg = "true";
defparam \entry_0[46] .power_up = "low";

cycloneive_lcell_comb \rd_address~0 (
	.dataa(\rd_address~q ),
	.datab(pending),
	.datac(gnd),
	.datad(f_pop),
	.cin(gnd),
	.combout(\rd_address~0_combout ),
	.cout());
defparam \rd_address~0 .lut_mask = 16'h9966;
defparam \rd_address~0 .sum_lutc_input = "datac";

dffeas rd_address(
	.clk(clk),
	.d(\rd_address~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_address~q ),
	.prn(vcc));
defparam rd_address.is_wysiwyg = "true";
defparam rd_address.power_up = "low";

dffeas \entry_1[61] (
	.clk(clk),
	.d(m0_write),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[61]~q ),
	.prn(vcc));
defparam \entry_1[61] .is_wysiwyg = "true";
defparam \entry_1[61] .power_up = "low";

dffeas \entry_0[61] (
	.clk(clk),
	.d(m0_write),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[61]~q ),
	.prn(vcc));
defparam \entry_0[61] .is_wysiwyg = "true";
defparam \entry_0[61] .power_up = "low";

dffeas \entry_1[60] (
	.clk(clk),
	.d(src_data_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[60]~q ),
	.prn(vcc));
defparam \entry_1[60] .is_wysiwyg = "true";
defparam \entry_1[60] .power_up = "low";

dffeas \entry_0[60] (
	.clk(clk),
	.d(src_data_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[60]~q ),
	.prn(vcc));
defparam \entry_0[60] .is_wysiwyg = "true";
defparam \entry_0[60] .power_up = "low";

dffeas \entry_1[47] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[47]~q ),
	.prn(vcc));
defparam \entry_1[47] .is_wysiwyg = "true";
defparam \entry_1[47] .power_up = "low";

dffeas \entry_0[47] (
	.clk(clk),
	.d(src_data_49),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[47]~q ),
	.prn(vcc));
defparam \entry_0[47] .is_wysiwyg = "true";
defparam \entry_0[47] .power_up = "low";

dffeas \entry_1[49] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[49]~q ),
	.prn(vcc));
defparam \entry_1[49] .is_wysiwyg = "true";
defparam \entry_1[49] .power_up = "low";

dffeas \entry_0[49] (
	.clk(clk),
	.d(src_data_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[49]~q ),
	.prn(vcc));
defparam \entry_0[49] .is_wysiwyg = "true";
defparam \entry_0[49] .power_up = "low";

dffeas \entry_1[48] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[48]~q ),
	.prn(vcc));
defparam \entry_1[48] .is_wysiwyg = "true";
defparam \entry_1[48] .power_up = "low";

dffeas \entry_0[48] (
	.clk(clk),
	.d(src_data_50),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[48]~q ),
	.prn(vcc));
defparam \entry_0[48] .is_wysiwyg = "true";
defparam \entry_0[48] .power_up = "low";

dffeas \entry_1[51] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[51]~q ),
	.prn(vcc));
defparam \entry_1[51] .is_wysiwyg = "true";
defparam \entry_1[51] .power_up = "low";

dffeas \entry_0[51] (
	.clk(clk),
	.d(src_data_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[51]~q ),
	.prn(vcc));
defparam \entry_0[51] .is_wysiwyg = "true";
defparam \entry_0[51] .power_up = "low";

dffeas \entry_1[50] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[50]~q ),
	.prn(vcc));
defparam \entry_1[50] .is_wysiwyg = "true";
defparam \entry_1[50] .power_up = "low";

dffeas \entry_0[50] (
	.clk(clk),
	.d(src_data_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[50]~q ),
	.prn(vcc));
defparam \entry_0[50] .is_wysiwyg = "true";
defparam \entry_0[50] .power_up = "low";

dffeas \entry_1[53] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[53]~q ),
	.prn(vcc));
defparam \entry_1[53] .is_wysiwyg = "true";
defparam \entry_1[53] .power_up = "low";

dffeas \entry_0[53] (
	.clk(clk),
	.d(src_data_55),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[53]~q ),
	.prn(vcc));
defparam \entry_0[53] .is_wysiwyg = "true";
defparam \entry_0[53] .power_up = "low";

dffeas \entry_1[52] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[52]~q ),
	.prn(vcc));
defparam \entry_1[52] .is_wysiwyg = "true";
defparam \entry_1[52] .power_up = "low";

dffeas \entry_0[52] (
	.clk(clk),
	.d(src_data_54),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[52]~q ),
	.prn(vcc));
defparam \entry_0[52] .is_wysiwyg = "true";
defparam \entry_0[52] .power_up = "low";

dffeas \entry_1[55] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[55]~q ),
	.prn(vcc));
defparam \entry_1[55] .is_wysiwyg = "true";
defparam \entry_1[55] .power_up = "low";

dffeas \entry_0[55] (
	.clk(clk),
	.d(src_data_57),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[55]~q ),
	.prn(vcc));
defparam \entry_0[55] .is_wysiwyg = "true";
defparam \entry_0[55] .power_up = "low";

dffeas \entry_1[54] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[54]~q ),
	.prn(vcc));
defparam \entry_1[54] .is_wysiwyg = "true";
defparam \entry_1[54] .power_up = "low";

dffeas \entry_0[54] (
	.clk(clk),
	.d(src_data_56),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[54]~q ),
	.prn(vcc));
defparam \entry_0[54] .is_wysiwyg = "true";
defparam \entry_0[54] .power_up = "low";

dffeas \entry_1[57] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[57]~q ),
	.prn(vcc));
defparam \entry_1[57] .is_wysiwyg = "true";
defparam \entry_1[57] .power_up = "low";

dffeas \entry_0[57] (
	.clk(clk),
	.d(src_data_59),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[57]~q ),
	.prn(vcc));
defparam \entry_0[57] .is_wysiwyg = "true";
defparam \entry_0[57] .power_up = "low";

dffeas \entry_1[56] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[56]~q ),
	.prn(vcc));
defparam \entry_1[56] .is_wysiwyg = "true";
defparam \entry_1[56] .power_up = "low";

dffeas \entry_0[56] (
	.clk(clk),
	.d(src_data_58),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[56]~q ),
	.prn(vcc));
defparam \entry_0[56] .is_wysiwyg = "true";
defparam \entry_0[56] .power_up = "low";

dffeas \entry_1[59] (
	.clk(clk),
	.d(src_data_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[59]~q ),
	.prn(vcc));
defparam \entry_1[59] .is_wysiwyg = "true";
defparam \entry_1[59] .power_up = "low";

dffeas \entry_0[59] (
	.clk(clk),
	.d(src_data_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[59]~q ),
	.prn(vcc));
defparam \entry_0[59] .is_wysiwyg = "true";
defparam \entry_0[59] .power_up = "low";

dffeas \entry_1[58] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[58]~q ),
	.prn(vcc));
defparam \entry_1[58] .is_wysiwyg = "true";
defparam \entry_1[58] .power_up = "low";

dffeas \entry_0[58] (
	.clk(clk),
	.d(src_data_60),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[58]~q ),
	.prn(vcc));
defparam \entry_0[58] .is_wysiwyg = "true";
defparam \entry_0[58] .power_up = "low";

dffeas \entry_1[36] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[36]~q ),
	.prn(vcc));
defparam \entry_1[36] .is_wysiwyg = "true";
defparam \entry_1[36] .power_up = "low";

dffeas \entry_0[36] (
	.clk(clk),
	.d(src_data_38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[36]~q ),
	.prn(vcc));
defparam \entry_0[36] .is_wysiwyg = "true";
defparam \entry_0[36] .power_up = "low";

dffeas \entry_1[37] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[37]~q ),
	.prn(vcc));
defparam \entry_1[37] .is_wysiwyg = "true";
defparam \entry_1[37] .power_up = "low";

dffeas \entry_0[37] (
	.clk(clk),
	.d(src_data_39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[37]~q ),
	.prn(vcc));
defparam \entry_0[37] .is_wysiwyg = "true";
defparam \entry_0[37] .power_up = "low";

dffeas \entry_1[38] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[38]~q ),
	.prn(vcc));
defparam \entry_1[38] .is_wysiwyg = "true";
defparam \entry_1[38] .power_up = "low";

dffeas \entry_0[38] (
	.clk(clk),
	.d(src_data_40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[38]~q ),
	.prn(vcc));
defparam \entry_0[38] .is_wysiwyg = "true";
defparam \entry_0[38] .power_up = "low";

dffeas \entry_1[39] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[39]~q ),
	.prn(vcc));
defparam \entry_1[39] .is_wysiwyg = "true";
defparam \entry_1[39] .power_up = "low";

dffeas \entry_0[39] (
	.clk(clk),
	.d(src_data_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[39]~q ),
	.prn(vcc));
defparam \entry_0[39] .is_wysiwyg = "true";
defparam \entry_0[39] .power_up = "low";

dffeas \entry_1[40] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[40]~q ),
	.prn(vcc));
defparam \entry_1[40] .is_wysiwyg = "true";
defparam \entry_1[40] .power_up = "low";

dffeas \entry_0[40] (
	.clk(clk),
	.d(src_data_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[40]~q ),
	.prn(vcc));
defparam \entry_0[40] .is_wysiwyg = "true";
defparam \entry_0[40] .power_up = "low";

dffeas \entry_1[41] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[41]~q ),
	.prn(vcc));
defparam \entry_1[41] .is_wysiwyg = "true";
defparam \entry_1[41] .power_up = "low";

dffeas \entry_0[41] (
	.clk(clk),
	.d(src_data_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[41]~q ),
	.prn(vcc));
defparam \entry_0[41] .is_wysiwyg = "true";
defparam \entry_0[41] .power_up = "low";

dffeas \entry_1[42] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[42]~q ),
	.prn(vcc));
defparam \entry_1[42] .is_wysiwyg = "true";
defparam \entry_1[42] .power_up = "low";

dffeas \entry_0[42] (
	.clk(clk),
	.d(src_data_44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[42]~q ),
	.prn(vcc));
defparam \entry_0[42] .is_wysiwyg = "true";
defparam \entry_0[42] .power_up = "low";

dffeas \entry_1[43] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[43]~q ),
	.prn(vcc));
defparam \entry_1[43] .is_wysiwyg = "true";
defparam \entry_1[43] .power_up = "low";

dffeas \entry_0[43] (
	.clk(clk),
	.d(src_data_45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[43]~q ),
	.prn(vcc));
defparam \entry_0[43] .is_wysiwyg = "true";
defparam \entry_0[43] .power_up = "low";

dffeas \entry_1[44] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[44]~q ),
	.prn(vcc));
defparam \entry_1[44] .is_wysiwyg = "true";
defparam \entry_1[44] .power_up = "low";

dffeas \entry_0[44] (
	.clk(clk),
	.d(src_data_46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[44]~q ),
	.prn(vcc));
defparam \entry_0[44] .is_wysiwyg = "true";
defparam \entry_0[44] .power_up = "low";

dffeas \entry_1[45] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[45]~q ),
	.prn(vcc));
defparam \entry_1[45] .is_wysiwyg = "true";
defparam \entry_1[45] .power_up = "low";

dffeas \entry_0[45] (
	.clk(clk),
	.d(src_data_47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[45]~q ),
	.prn(vcc));
defparam \entry_0[45] .is_wysiwyg = "true";
defparam \entry_0[45] .power_up = "low";

dffeas \entry_1[32] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[32]~q ),
	.prn(vcc));
defparam \entry_1[32] .is_wysiwyg = "true";
defparam \entry_1[32] .power_up = "low";

dffeas \entry_0[32] (
	.clk(clk),
	.d(comb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[32]~q ),
	.prn(vcc));
defparam \entry_0[32] .is_wysiwyg = "true";
defparam \entry_0[32] .power_up = "low";

dffeas \entry_1[33] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[33]~q ),
	.prn(vcc));
defparam \entry_1[33] .is_wysiwyg = "true";
defparam \entry_1[33] .power_up = "low";

dffeas \entry_0[33] (
	.clk(clk),
	.d(comb1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[33]~q ),
	.prn(vcc));
defparam \entry_0[33] .is_wysiwyg = "true";
defparam \entry_0[33] .power_up = "low";

dffeas \entry_1[34] (
	.clk(clk),
	.d(comb2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[34]~q ),
	.prn(vcc));
defparam \entry_1[34] .is_wysiwyg = "true";
defparam \entry_1[34] .power_up = "low";

dffeas \entry_0[34] (
	.clk(clk),
	.d(comb2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[34]~q ),
	.prn(vcc));
defparam \entry_0[34] .is_wysiwyg = "true";
defparam \entry_0[34] .power_up = "low";

dffeas \entry_1[35] (
	.clk(clk),
	.d(comb3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[35]~q ),
	.prn(vcc));
defparam \entry_1[35] .is_wysiwyg = "true";
defparam \entry_1[35] .power_up = "low";

dffeas \entry_0[35] (
	.clk(clk),
	.d(comb3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[35]~q ),
	.prn(vcc));
defparam \entry_0[35] .is_wysiwyg = "true";
defparam \entry_0[35] .power_up = "low";

dffeas \entry_1[0] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[0]~q ),
	.prn(vcc));
defparam \entry_1[0] .is_wysiwyg = "true";
defparam \entry_1[0] .power_up = "low";

dffeas \entry_0[0] (
	.clk(clk),
	.d(src_payload1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[0]~q ),
	.prn(vcc));
defparam \entry_0[0] .is_wysiwyg = "true";
defparam \entry_0[0] .power_up = "low";

dffeas \entry_1[1] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[1]~q ),
	.prn(vcc));
defparam \entry_1[1] .is_wysiwyg = "true";
defparam \entry_1[1] .power_up = "low";

dffeas \entry_0[1] (
	.clk(clk),
	.d(src_payload2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[1]~q ),
	.prn(vcc));
defparam \entry_0[1] .is_wysiwyg = "true";
defparam \entry_0[1] .power_up = "low";

dffeas \entry_1[2] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[2]~q ),
	.prn(vcc));
defparam \entry_1[2] .is_wysiwyg = "true";
defparam \entry_1[2] .power_up = "low";

dffeas \entry_0[2] (
	.clk(clk),
	.d(src_payload3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[2]~q ),
	.prn(vcc));
defparam \entry_0[2] .is_wysiwyg = "true";
defparam \entry_0[2] .power_up = "low";

dffeas \entry_1[3] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[3]~q ),
	.prn(vcc));
defparam \entry_1[3] .is_wysiwyg = "true";
defparam \entry_1[3] .power_up = "low";

dffeas \entry_0[3] (
	.clk(clk),
	.d(src_payload4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[3]~q ),
	.prn(vcc));
defparam \entry_0[3] .is_wysiwyg = "true";
defparam \entry_0[3] .power_up = "low";

dffeas \entry_1[4] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[4]~q ),
	.prn(vcc));
defparam \entry_1[4] .is_wysiwyg = "true";
defparam \entry_1[4] .power_up = "low";

dffeas \entry_0[4] (
	.clk(clk),
	.d(src_payload5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[4]~q ),
	.prn(vcc));
defparam \entry_0[4] .is_wysiwyg = "true";
defparam \entry_0[4] .power_up = "low";

dffeas \entry_1[5] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[5]~q ),
	.prn(vcc));
defparam \entry_1[5] .is_wysiwyg = "true";
defparam \entry_1[5] .power_up = "low";

dffeas \entry_0[5] (
	.clk(clk),
	.d(src_payload6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[5]~q ),
	.prn(vcc));
defparam \entry_0[5] .is_wysiwyg = "true";
defparam \entry_0[5] .power_up = "low";

dffeas \entry_1[6] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[6]~q ),
	.prn(vcc));
defparam \entry_1[6] .is_wysiwyg = "true";
defparam \entry_1[6] .power_up = "low";

dffeas \entry_0[6] (
	.clk(clk),
	.d(src_payload7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[6]~q ),
	.prn(vcc));
defparam \entry_0[6] .is_wysiwyg = "true";
defparam \entry_0[6] .power_up = "low";

dffeas \entry_1[7] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[7]~q ),
	.prn(vcc));
defparam \entry_1[7] .is_wysiwyg = "true";
defparam \entry_1[7] .power_up = "low";

dffeas \entry_0[7] (
	.clk(clk),
	.d(src_payload8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[7]~q ),
	.prn(vcc));
defparam \entry_0[7] .is_wysiwyg = "true";
defparam \entry_0[7] .power_up = "low";

dffeas \entry_1[8] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[8]~q ),
	.prn(vcc));
defparam \entry_1[8] .is_wysiwyg = "true";
defparam \entry_1[8] .power_up = "low";

dffeas \entry_0[8] (
	.clk(clk),
	.d(src_payload9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[8]~q ),
	.prn(vcc));
defparam \entry_0[8] .is_wysiwyg = "true";
defparam \entry_0[8] .power_up = "low";

dffeas \entry_1[9] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[9]~q ),
	.prn(vcc));
defparam \entry_1[9] .is_wysiwyg = "true";
defparam \entry_1[9] .power_up = "low";

dffeas \entry_0[9] (
	.clk(clk),
	.d(src_payload10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[9]~q ),
	.prn(vcc));
defparam \entry_0[9] .is_wysiwyg = "true";
defparam \entry_0[9] .power_up = "low";

dffeas \entry_1[10] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[10]~q ),
	.prn(vcc));
defparam \entry_1[10] .is_wysiwyg = "true";
defparam \entry_1[10] .power_up = "low";

dffeas \entry_0[10] (
	.clk(clk),
	.d(src_payload11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[10]~q ),
	.prn(vcc));
defparam \entry_0[10] .is_wysiwyg = "true";
defparam \entry_0[10] .power_up = "low";

dffeas \entry_1[11] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[11]~q ),
	.prn(vcc));
defparam \entry_1[11] .is_wysiwyg = "true";
defparam \entry_1[11] .power_up = "low";

dffeas \entry_0[11] (
	.clk(clk),
	.d(src_payload12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[11]~q ),
	.prn(vcc));
defparam \entry_0[11] .is_wysiwyg = "true";
defparam \entry_0[11] .power_up = "low";

dffeas \entry_1[12] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[12]~q ),
	.prn(vcc));
defparam \entry_1[12] .is_wysiwyg = "true";
defparam \entry_1[12] .power_up = "low";

dffeas \entry_0[12] (
	.clk(clk),
	.d(src_payload13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[12]~q ),
	.prn(vcc));
defparam \entry_0[12] .is_wysiwyg = "true";
defparam \entry_0[12] .power_up = "low";

dffeas \entry_1[13] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[13]~q ),
	.prn(vcc));
defparam \entry_1[13] .is_wysiwyg = "true";
defparam \entry_1[13] .power_up = "low";

dffeas \entry_0[13] (
	.clk(clk),
	.d(src_payload14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[13]~q ),
	.prn(vcc));
defparam \entry_0[13] .is_wysiwyg = "true";
defparam \entry_0[13] .power_up = "low";

dffeas \entry_1[14] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[14]~q ),
	.prn(vcc));
defparam \entry_1[14] .is_wysiwyg = "true";
defparam \entry_1[14] .power_up = "low";

dffeas \entry_0[14] (
	.clk(clk),
	.d(src_payload15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[14]~q ),
	.prn(vcc));
defparam \entry_0[14] .is_wysiwyg = "true";
defparam \entry_0[14] .power_up = "low";

dffeas \entry_1[15] (
	.clk(clk),
	.d(src_payload16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[15]~q ),
	.prn(vcc));
defparam \entry_1[15] .is_wysiwyg = "true";
defparam \entry_1[15] .power_up = "low";

dffeas \entry_0[15] (
	.clk(clk),
	.d(src_payload16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[15]~q ),
	.prn(vcc));
defparam \entry_0[15] .is_wysiwyg = "true";
defparam \entry_0[15] .power_up = "low";

dffeas \entry_1[16] (
	.clk(clk),
	.d(src_payload17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[16]~q ),
	.prn(vcc));
defparam \entry_1[16] .is_wysiwyg = "true";
defparam \entry_1[16] .power_up = "low";

dffeas \entry_0[16] (
	.clk(clk),
	.d(src_payload17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[16]~q ),
	.prn(vcc));
defparam \entry_0[16] .is_wysiwyg = "true";
defparam \entry_0[16] .power_up = "low";

dffeas \entry_1[17] (
	.clk(clk),
	.d(src_payload18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[17]~q ),
	.prn(vcc));
defparam \entry_1[17] .is_wysiwyg = "true";
defparam \entry_1[17] .power_up = "low";

dffeas \entry_0[17] (
	.clk(clk),
	.d(src_payload18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[17]~q ),
	.prn(vcc));
defparam \entry_0[17] .is_wysiwyg = "true";
defparam \entry_0[17] .power_up = "low";

dffeas \entry_1[18] (
	.clk(clk),
	.d(src_payload19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[18]~q ),
	.prn(vcc));
defparam \entry_1[18] .is_wysiwyg = "true";
defparam \entry_1[18] .power_up = "low";

dffeas \entry_0[18] (
	.clk(clk),
	.d(src_payload19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[18]~q ),
	.prn(vcc));
defparam \entry_0[18] .is_wysiwyg = "true";
defparam \entry_0[18] .power_up = "low";

dffeas \entry_1[19] (
	.clk(clk),
	.d(src_payload20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[19]~q ),
	.prn(vcc));
defparam \entry_1[19] .is_wysiwyg = "true";
defparam \entry_1[19] .power_up = "low";

dffeas \entry_0[19] (
	.clk(clk),
	.d(src_payload20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[19]~q ),
	.prn(vcc));
defparam \entry_0[19] .is_wysiwyg = "true";
defparam \entry_0[19] .power_up = "low";

dffeas \entry_1[20] (
	.clk(clk),
	.d(src_payload21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[20]~q ),
	.prn(vcc));
defparam \entry_1[20] .is_wysiwyg = "true";
defparam \entry_1[20] .power_up = "low";

dffeas \entry_0[20] (
	.clk(clk),
	.d(src_payload21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[20]~q ),
	.prn(vcc));
defparam \entry_0[20] .is_wysiwyg = "true";
defparam \entry_0[20] .power_up = "low";

dffeas \entry_1[21] (
	.clk(clk),
	.d(src_payload22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[21]~q ),
	.prn(vcc));
defparam \entry_1[21] .is_wysiwyg = "true";
defparam \entry_1[21] .power_up = "low";

dffeas \entry_0[21] (
	.clk(clk),
	.d(src_payload22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[21]~q ),
	.prn(vcc));
defparam \entry_0[21] .is_wysiwyg = "true";
defparam \entry_0[21] .power_up = "low";

dffeas \entry_1[22] (
	.clk(clk),
	.d(src_payload23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[22]~q ),
	.prn(vcc));
defparam \entry_1[22] .is_wysiwyg = "true";
defparam \entry_1[22] .power_up = "low";

dffeas \entry_0[22] (
	.clk(clk),
	.d(src_payload23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[22]~q ),
	.prn(vcc));
defparam \entry_0[22] .is_wysiwyg = "true";
defparam \entry_0[22] .power_up = "low";

dffeas \entry_1[23] (
	.clk(clk),
	.d(src_payload24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[23]~q ),
	.prn(vcc));
defparam \entry_1[23] .is_wysiwyg = "true";
defparam \entry_1[23] .power_up = "low";

dffeas \entry_0[23] (
	.clk(clk),
	.d(src_payload24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[23]~q ),
	.prn(vcc));
defparam \entry_0[23] .is_wysiwyg = "true";
defparam \entry_0[23] .power_up = "low";

dffeas \entry_1[24] (
	.clk(clk),
	.d(src_payload25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[24]~q ),
	.prn(vcc));
defparam \entry_1[24] .is_wysiwyg = "true";
defparam \entry_1[24] .power_up = "low";

dffeas \entry_0[24] (
	.clk(clk),
	.d(src_payload25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[24]~q ),
	.prn(vcc));
defparam \entry_0[24] .is_wysiwyg = "true";
defparam \entry_0[24] .power_up = "low";

dffeas \entry_1[25] (
	.clk(clk),
	.d(src_payload26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[25]~q ),
	.prn(vcc));
defparam \entry_1[25] .is_wysiwyg = "true";
defparam \entry_1[25] .power_up = "low";

dffeas \entry_0[25] (
	.clk(clk),
	.d(src_payload26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[25]~q ),
	.prn(vcc));
defparam \entry_0[25] .is_wysiwyg = "true";
defparam \entry_0[25] .power_up = "low";

dffeas \entry_1[26] (
	.clk(clk),
	.d(src_payload27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[26]~q ),
	.prn(vcc));
defparam \entry_1[26] .is_wysiwyg = "true";
defparam \entry_1[26] .power_up = "low";

dffeas \entry_0[26] (
	.clk(clk),
	.d(src_payload27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[26]~q ),
	.prn(vcc));
defparam \entry_0[26] .is_wysiwyg = "true";
defparam \entry_0[26] .power_up = "low";

dffeas \entry_1[27] (
	.clk(clk),
	.d(src_payload28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[27]~q ),
	.prn(vcc));
defparam \entry_1[27] .is_wysiwyg = "true";
defparam \entry_1[27] .power_up = "low";

dffeas \entry_0[27] (
	.clk(clk),
	.d(src_payload28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[27]~q ),
	.prn(vcc));
defparam \entry_0[27] .is_wysiwyg = "true";
defparam \entry_0[27] .power_up = "low";

dffeas \entry_1[28] (
	.clk(clk),
	.d(src_payload29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[28]~q ),
	.prn(vcc));
defparam \entry_1[28] .is_wysiwyg = "true";
defparam \entry_1[28] .power_up = "low";

dffeas \entry_0[28] (
	.clk(clk),
	.d(src_payload29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[28]~q ),
	.prn(vcc));
defparam \entry_0[28] .is_wysiwyg = "true";
defparam \entry_0[28] .power_up = "low";

dffeas \entry_1[29] (
	.clk(clk),
	.d(src_payload30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[29]~q ),
	.prn(vcc));
defparam \entry_1[29] .is_wysiwyg = "true";
defparam \entry_1[29] .power_up = "low";

dffeas \entry_0[29] (
	.clk(clk),
	.d(src_payload30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[29]~q ),
	.prn(vcc));
defparam \entry_0[29] .is_wysiwyg = "true";
defparam \entry_0[29] .power_up = "low";

dffeas \entry_1[30] (
	.clk(clk),
	.d(src_payload31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[30]~q ),
	.prn(vcc));
defparam \entry_1[30] .is_wysiwyg = "true";
defparam \entry_1[30] .power_up = "low";

dffeas \entry_0[30] (
	.clk(clk),
	.d(src_payload31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[30]~q ),
	.prn(vcc));
defparam \entry_0[30] .is_wysiwyg = "true";
defparam \entry_0[30] .power_up = "low";

dffeas \entry_1[31] (
	.clk(clk),
	.d(src_payload32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_1[61]~0_combout ),
	.q(\entry_1[31]~q ),
	.prn(vcc));
defparam \entry_1[31] .is_wysiwyg = "true";
defparam \entry_1[31] .power_up = "low";

dffeas \entry_0[31] (
	.clk(clk),
	.d(src_payload32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entry_0[61]~0_combout ),
	.q(\entry_0[31]~q ),
	.prn(vcc));
defparam \entry_0[31] .is_wysiwyg = "true";
defparam \entry_0[31] .power_up = "low";

endmodule

module final_project_soc_final_project_soc_sdram_pll (
	wire_pll7_clk_0,
	wire_pll7_clk_1,
	locked,
	d_writedata_0,
	reset,
	d_writedata_1,
	mem_used_1,
	WideOr1,
	src_data_38,
	mem,
	src_data_39,
	mem1,
	readdata_0,
	readdata_1,
	clk_clk,
	unused_sdram_areset_conduit_export)/* synthesis synthesis_greybox=1 */;
output 	wire_pll7_clk_0;
output 	wire_pll7_clk_1;
output 	locked;
input 	d_writedata_0;
input 	reset;
input 	d_writedata_1;
input 	mem_used_1;
input 	WideOr1;
input 	src_data_38;
input 	mem;
input 	src_data_39;
input 	mem1;
output 	readdata_0;
output 	readdata_1;
input 	clk_clk;
input 	unused_sdram_areset_conduit_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \comb~0_combout ;
wire \stdsync2|dffpipe3|dffe6a[0]~q ;
wire \readdata[0]~0_combout ;
wire \w_reset~0_combout ;
wire \w_reset~1_combout ;
wire \prev_reset~q ;
wire \pfdena_reg~0_combout ;
wire \pfdena_reg~q ;


final_project_soc_final_project_soc_sdram_pll_altpll_fua2 sd1(
	.clk({clk_unconnected_wire_4,clk_unconnected_wire_3,clk_unconnected_wire_2,wire_pll7_clk_1,wire_pll7_clk_0}),
	.locked1(locked),
	.areset(\comb~0_combout ),
	.inclk({gnd,clk_clk}));

final_project_soc_final_project_soc_sdram_pll_stdsync_sv6 stdsync2(
	.locked(locked),
	.r_sync_rst(reset),
	.dffe6a_0(\stdsync2|dffpipe3|dffe6a[0]~q ),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \comb~0 (
	.dataa(unused_sdram_areset_conduit_export),
	.datab(\prev_reset~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'hEEEE;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~1 (
	.dataa(\readdata[0]~0_combout ),
	.datab(\prev_reset~q ),
	.datac(\stdsync2|dffpipe3|dffe6a[0]~q ),
	.datad(src_data_38),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0]~1 .lut_mask = 16'hFAFC;
defparam \readdata[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1]~2 (
	.dataa(\readdata[0]~0_combout ),
	.datab(gnd),
	.datac(src_data_38),
	.datad(\pfdena_reg~q ),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1]~2 .lut_mask = 16'hAFFF;
defparam \readdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0]~0 (
	.dataa(WideOr1),
	.datab(mem1),
	.datac(mem_used_1),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\readdata[0]~0_combout ),
	.cout());
defparam \readdata[0]~0 .lut_mask = 16'hEFFF;
defparam \readdata[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \w_reset~0 (
	.dataa(WideOr1),
	.datab(src_data_38),
	.datac(mem),
	.datad(src_data_39),
	.cin(gnd),
	.combout(\w_reset~0_combout ),
	.cout());
defparam \w_reset~0 .lut_mask = 16'hFEFF;
defparam \w_reset~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \w_reset~1 (
	.dataa(d_writedata_0),
	.datab(\w_reset~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\w_reset~1_combout ),
	.cout());
defparam \w_reset~1 .lut_mask = 16'hEEEE;
defparam \w_reset~1 .sum_lutc_input = "datac";

dffeas prev_reset(
	.clk(clk_clk),
	.d(\w_reset~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prev_reset~q ),
	.prn(vcc));
defparam prev_reset.is_wysiwyg = "true";
defparam prev_reset.power_up = "low";

cycloneive_lcell_comb \pfdena_reg~0 (
	.dataa(d_writedata_1),
	.datab(\w_reset~0_combout ),
	.datac(gnd),
	.datad(\pfdena_reg~q ),
	.cin(gnd),
	.combout(\pfdena_reg~0_combout ),
	.cout());
defparam \pfdena_reg~0 .lut_mask = 16'hDD11;
defparam \pfdena_reg~0 .sum_lutc_input = "datac";

dffeas pfdena_reg(
	.clk(clk_clk),
	.d(\pfdena_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pfdena_reg~q ),
	.prn(vcc));
defparam pfdena_reg.is_wysiwyg = "true";
defparam pfdena_reg.power_up = "low";

endmodule

module final_project_soc_final_project_soc_sdram_pll_altpll_fua2 (
	clk,
	locked1,
	areset,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	[4:0] clk;
output 	locked1;
input 	areset;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wire_pll7_clk[2] ;
wire \wire_pll7_clk[3] ;
wire \wire_pll7_clk[4] ;
wire wire_pll7_locked;
wire wire_pll7_fbout;
wire \pll_lock_sync~q ;

wire [4:0] pll7_CLK_bus;

assign clk[0] = pll7_CLK_bus[0];
assign clk[1] = pll7_CLK_bus[1];
assign \wire_pll7_clk[2]  = pll7_CLK_bus[2];
assign \wire_pll7_clk[3]  = pll7_CLK_bus[3];
assign \wire_pll7_clk[4]  = pll7_CLK_bus[4];

cycloneive_pll pll7(
	.areset(areset),
	.pfdena(vcc),
	.fbin(wire_pll7_fbout),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scandata(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect(3'b000),
	.phasedone(),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(wire_pll7_locked),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(wire_pll7_fbout),
	.clk(pll7_CLK_bus),
	.clkbad());
defparam pll7.auto_settings = "false";
defparam pll7.bandwidth_type = "auto";
defparam pll7.c0_high = 10;
defparam pll7.c0_initial = 4;
defparam pll7.c0_low = 10;
defparam pll7.c0_mode = "even";
defparam pll7.c0_ph = 0;
defparam pll7.c1_high = 10;
defparam pll7.c1_initial = 1;
defparam pll7.c1_low = 10;
defparam pll7.c1_mode = "even";
defparam pll7.c1_ph = 0;
defparam pll7.c1_use_casc_in = "off";
defparam pll7.c2_high = 1;
defparam pll7.c2_initial = 1;
defparam pll7.c2_low = 1;
defparam pll7.c2_mode = "bypass";
defparam pll7.c2_ph = 0;
defparam pll7.c2_use_casc_in = "off";
defparam pll7.c3_high = 1;
defparam pll7.c3_initial = 1;
defparam pll7.c3_low = 1;
defparam pll7.c3_mode = "bypass";
defparam pll7.c3_ph = 0;
defparam pll7.c3_use_casc_in = "off";
defparam pll7.c4_high = 1;
defparam pll7.c4_initial = 1;
defparam pll7.c4_low = 1;
defparam pll7.c4_mode = "bypass";
defparam pll7.c4_ph = 0;
defparam pll7.c4_use_casc_in = "off";
defparam pll7.charge_pump_current_bits = 2;
defparam pll7.clk0_counter = "c0";
defparam pll7.clk0_divide_by = 1;
defparam pll7.clk0_duty_cycle = 50;
defparam pll7.clk0_multiply_by = 1;
defparam pll7.clk0_phase_shift = "0";
defparam pll7.clk1_counter = "c1";
defparam pll7.clk1_divide_by = 1;
defparam pll7.clk1_duty_cycle = 50;
defparam pll7.clk1_multiply_by = 1;
defparam pll7.clk1_phase_shift = "-3000";
defparam pll7.clk2_counter = "unused";
defparam pll7.clk2_divide_by = 0;
defparam pll7.clk2_duty_cycle = 50;
defparam pll7.clk2_multiply_by = 0;
defparam pll7.clk2_phase_shift = "0";
defparam pll7.clk3_counter = "unused";
defparam pll7.clk3_divide_by = 0;
defparam pll7.clk3_duty_cycle = 50;
defparam pll7.clk3_multiply_by = 0;
defparam pll7.clk3_phase_shift = "0";
defparam pll7.clk4_counter = "unused";
defparam pll7.clk4_divide_by = 0;
defparam pll7.clk4_duty_cycle = 50;
defparam pll7.clk4_multiply_by = 0;
defparam pll7.clk4_phase_shift = "0";
defparam pll7.compensate_clock = "clock0";
defparam pll7.inclk0_input_frequency = 20000;
defparam pll7.inclk1_input_frequency = 0;
defparam pll7.loop_filter_c_bits = 2;
defparam pll7.loop_filter_r_bits = 1;
defparam pll7.m = 20;
defparam pll7.m_initial = 4;
defparam pll7.m_ph = 0;
defparam pll7.n = 1;
defparam pll7.operation_mode = "normal";
defparam pll7.pfd_max = 0;
defparam pll7.pfd_min = 0;
defparam pll7.self_reset_on_loss_lock = "off";
defparam pll7.simulation_type = "timing";
defparam pll7.switch_over_type = "auto";
defparam pll7.vco_center = 0;
defparam pll7.vco_divide_by = 0;
defparam pll7.vco_frequency_control = "auto";
defparam pll7.vco_max = 0;
defparam pll7.vco_min = 0;
defparam pll7.vco_multiply_by = 0;
defparam pll7.vco_phase_shift_step = 0;
defparam pll7.vco_post_scale = 1;

cycloneive_lcell_comb locked(
	.dataa(wire_pll7_locked),
	.datab(\pll_lock_sync~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(locked1),
	.cout());
defparam locked.lut_mask = 16'hEEEE;
defparam locked.sum_lutc_input = "datac";

dffeas pll_lock_sync(
	.clk(wire_pll7_locked),
	.d(vcc),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_lock_sync~q ),
	.prn(vcc));
defparam pll_lock_sync.is_wysiwyg = "true";
defparam pll_lock_sync.power_up = "low";

endmodule

module final_project_soc_final_project_soc_sdram_pll_stdsync_sv6 (
	locked,
	r_sync_rst,
	dffe6a_0,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	locked;
input 	r_sync_rst;
output 	dffe6a_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



final_project_soc_final_project_soc_sdram_pll_dffpipe_l2c dffpipe3(
	.d({locked}),
	.clrn(r_sync_rst),
	.dffe6a_0(dffe6a_0),
	.clock(clk_clk));

endmodule

module final_project_soc_final_project_soc_sdram_pll_dffpipe_l2c (
	d,
	clrn,
	dffe6a_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[0:0] d;
input 	clrn;
output 	dffe6a_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe4a[0]~q ;
wire \dffe5a[0]~q ;


dffeas \dffe6a[0] (
	.clk(clock),
	.d(\dffe5a[0]~q ),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe6a_0),
	.prn(vcc));
defparam \dffe6a[0] .is_wysiwyg = "true";
defparam \dffe6a[0] .power_up = "low";

dffeas \dffe4a[0] (
	.clk(clock),
	.d(d[0]),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe4a[0]~q ),
	.prn(vcc));
defparam \dffe4a[0] .is_wysiwyg = "true";
defparam \dffe4a[0] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock),
	.d(\dffe4a[0]~q ),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe5a[0]~q ),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

endmodule
